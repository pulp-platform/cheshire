/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module /scratch/zexifu/c910_pulp/merge_with_cyril/cheshire_with_c910/target/sim/src/dpi/bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 883;

    const logic [RomSize-1:0][63:0] mem = {
        64'h02faf080_00bebc20,
        64'h00001500_02000050,
        64'h00007700_00004069,
        64'h000087aa_01000048,
        64'h02faf080_00030d40,
        64'h622c4101_1494cf98,
        64'h4ce4fd95_0269b26a,
        64'h54524150_20494645,
        64'h00000000_00000005,
        64'h00000000_00000005,
        64'h00000000_00000002,
        64'h00000000_00000001,
        64'h00000000_00000001,
        64'hf2e0d6c4_baa89e8c,
        64'h62704654_2a380e1c,
        64'hc0d2e4f6_889aacbe,
        64'h50427466_180a3c2e,
        64'h9684b2a0_deccfae8,
        64'h06142230_4e5c6a78,
        64'ha4b68092_ecfec8da,
        64'h34261002_7c6e584a,
        64'h3a281e0c_72605644,
        64'haab88e9c_e2f0c6d4,
        64'h081a2c3e_40526476,
        64'h988abcae_d0c2f4e6,
        64'h5e4c7a68_16043220,
        64'hcedceaf8_8694a2b0,
        64'h6c7e485a_24360012,
        64'hfceed8ca_b4a69082,
        64'h70625446_382a1c0e,
        64'he0f2c4d6_a8ba8c9e,
        64'h42506674_0a182e3c,
        64'hd2c0f6e4_9a88beac,
        64'h14063022_5c4e786a,
        64'h8496a0b2_ccdee8fa,
        64'h26340210_6e7c4a58,
        64'hb6a49280_feecdac8,
        64'hb8aa9c8e_f0e2d4c6,
        64'h283a0c1e_60724456,
        64'h8a98aebc_c2d0e6f4,
        64'h1a083e2c_52407664,
        64'hdccef8ea_9486b0a2,
        64'h4c5e687a_04162032,
        64'heefccad8_a6b48290,
        64'h7e6c5a48_36241200,
        64'h1ef00ed1_3eb22e93,
        64'h5e744e55_7e366e17,
        64'h9ff88fd9_bfbaaf9b,
        64'hdf7ccf5d_ff3eef1f,
        64'h0cc11ce0_2c833ca2,
        64'h4c455c64_6c077c26,
        64'h8dc99de8_ad8bbdaa,
        64'hcd4ddd6c_ed0ffd2e,
        64'h3a922ab3_1ad00af1,
        64'h7a166a37_5a544a75,
        64'hbb9aabbb_9bd88bf9,
        64'hfb1eeb3f_db5ccb7d,
        64'h28a33882_08e118c0,
        64'h68277806_48655844,
        64'ha9abb98a_89e999c8,
        64'he92ff90e_c96dd94c,
        64'h56344615_76766657,
        64'h16b00691_36f226d3,
        64'hd73cc71d_f77ee75f,
        64'h97b88799_b7faa7db,
        64'h44055424_64477466,
        64'h048114a0_24c334e2,
        64'hc50dd52c_e54ff56e,
        64'h858995a8_a5cbb5ea,
        64'h72566277_52144235,
        64'h32d222f3_129002b1,
        64'hf35ee37f_d31cc33d,
        64'hb3daa3fb_939883b9,
        64'h60677046_40255004,
        64'h20e330c2_00a11080,
        64'he16ff14e_c12dd10c,
        64'ha1ebb1ca_81a99188,
        64'h8f789f59_af3abf1b,
        64'hcffcdfdd_efbeff9f,
        64'h0e701e51_2e323e13,
        64'h4ef45ed5_6eb67e97,
        64'h9d498d68_bd0bad2a,
        64'hddcdcdec_fd8fedae,
        64'h1c410c60_3c032c22,
        64'h5cc54ce4_7c876ca6,
        64'hab1abb3b_8b589b79,
        64'heb9efbbf_cbdcdbfd,
        64'h2a123a33_0a501a71,
        64'h6a967ab7_4ad45af5,
        64'hb92ba90a_99698948,
        64'hf9afe98e_d9edc9cc,
        64'h38232802_18610840,
        64'h78a76886_58e548c4,
        64'hc7bcd79d_e7fef7df,
        64'h87389719_a77ab75b,
        64'h46b45695_66f676d7,
        64'h06301611_26723653,
        64'hd58dc5ac_f5cfe5ee,
        64'h95098528_b54ba56a,
        64'h548544a4_74c764e6,
        64'h14010420_34432462,
        64'he3def3ff_c39cd3bd,
        64'ha35ab37b_83189339,
        64'h62d672f7_429452b5,
        64'h22523273_02101231,
        64'hf1efe1ce_d1adc18c,
        64'hb16ba14a_91298108,
        64'h70e760c6_50a54084,
        64'h30632042_10210000,
        64'h00000000_b595c085,
        64'h0513102c_cb98ffff,
        64'hf5170017_67137ee7,
        64'h87930100_17974b98,
        64'h7f878793_01001797,
        64'hc33c07f9_80470713,
        64'h01002717_df540695,
        64'h81270713_66c10100,
        64'h2717df14_06f98227,
        64'h0713001e_06b70100,
        64'h2717db54_06958327,
        64'h0713000f_06b70100,
        64'h2717db14_84070713,
        64'h02878693_01002717,
        64'h004107b7_d3981007,
        64'h67138527_87930100,
        64'h27975398_85c78793,
        64'h01002797_d3980017,
        64'h671386a7_87930100,
        64'h27975398_87478793,
        64'h01002797_d3980027,
        64'h67138827_87930100,
        64'h27975398_88c78793,
        64'h01002797_d3980807,
        64'h671389a7_87930100,
        64'h27975398_8a478793,
        64'h01002797_cb989b79,
        64'h8b078793_01002797,
        64'h4b988ba7_87930100,
        64'h2797f43e_8c478793,
        64'h01002797_bf913305,
        64'h0513102c_fffff517,
        64'ha93fe0ef_050502f5,
        64'h55332407_8793000f,
        64'h47b702f5_053315e0,
        64'h07939101_cb1c0204,
        64'h15138fa7_07130100,
        64'h37178fd9_20000737,
        64'h8ff9177d_e0000737,
        64'h4b9c9127_87930100,
        64'h3797cb98_80000737,
        64'h92078793_01003797,
        64'hf9552501_dc7fe0ef,
        64'he82e1028_46856662,
        64'h00011e23_cc3ef0f7,
        64'h8793000f_17b74d67,
        64'hb5830000_079784ef,
        64'hf0eff42a_fc3e4785,
        64'hf83e95a5_05130100,
        64'h3517c207_879300be,
        64'hc7b78082_61656946,
        64'h64e67406_70a6c0df,
        64'hf0efc0e5_0513080c,
        64'h00000517_b3ffe0ef,
        64'h050502f5_55332407,
        64'h8793000f_47b702f5,
        64'h05333e80_07939101,
        64'hc89c8fd9_0127f7b3,
        64'h02041513_20000737,
        64'h489ced1d_2501e51f,
        64'he0ef0808_66226582,
        64'h5692e539_2501e61f,
        64'he0ef6582_c03e5682,
        64'h67e2c89c_0127f7b3,
        64'h08086622_489c197d,
        64'he0000937_64c2e92d,
        64'h883ff0ef_08084601,
        64'h46854701_57c7b583,
        64'h00000797_e541899f,
        64'hf0ef0808_07a58593,
        64'h460d4681_470115a2,
        64'h0fd00593_fbf90281,
        64'h4783e15d_f56ff0ef,
        64'h08084601_10344701,
        64'h5a87b583_00000797,
        64'hed558cdf_f0ef0808,
        64'h85a64601_46814701,
        64'h07748493_14a20650,
        64'h04930291_0423ed69,
        64'h8ebff0ef_08084611,
        64'h46850705_07325da7,
        64'hb5830aa0_17370000,
        64'h07970e05_1c63909f,
        64'hf0ef0808_04058593,
        64'h46014685_470515a2,
        64'h09500593_10051963,
        64'h2501ef0f_f0effc3e,
        64'hd44ae482_e082f802,
        64'h08081030_46850500,
        64'h0793f402_5582cb1c,
        64'haa870713_01003717,
        64'h8fd92000_07378ff9,
        64'h177de000_07374b9c,
        64'hac078793_01003797,
        64'hcb988000_0737ace7,
        64'h87930100_37971605,
        64'h12632501_f77fe0ef,
        64'h08086622_65825692,
        64'h16051b63_2501f89f,
        64'he0efe402_e02e0808,
        64'h46014681_66c7b583,
        64'h00000797_a04ff0ef,
        64'hd24ad002_e82aec3e,
        64'hb1450513_60078793,
        64'h01003517_016e37b7,
        64'hb7096165_694664e6,
        64'h70a67406_00f48863,
        64'h478526f4_8563478d,
        64'h0007049b_1d270b63,
        64'h24014909_eca6f486,
        64'he8ca43e0_f0a2b507,
        64'h87937159_00fff797,
        64'h43b8b5a7_879300ff,
        64'hf7978b2f_f06ffae7,
        64'h98e3b6a7_c7830100,
        64'h1797dfcd_8b850147,
        64'hc783b7a7_87930100,
        64'h1797c3bf_e06f8d5d,
        64'h93811782_1502b8e7,
        64'ha78300ff_f79743c8,
        64'hb9878793_00fff797,
        64'h0007a423_ba478793,
        64'h00fff797_c7958b89,
        64'h479cbb27_879300ff,
        64'hf7974719_0ff0000f,
        64'h00e78823_02000713,
        64'hbc878793_01001797,
        64'h00e78423_fc700713,
        64'hbd878793_01001797,
        64'h00e78623_470dbe67,
        64'h87930100_17970007,
        64'h8223bf27_87930100,
        64'h1797bee7_8e23476d,
        64'h01001797_00e78623,
        64'hf8000713_c0c78793,
        64'h01001797_00078223,
        64'hc1878793_01001797,
        64'hb795f4f7_1fe37722,
        64'h7907b783_00000797,
        64'hce9fe06f_6165c385,
        64'h0513c7d8_0dfff517,
        64'hc5278793_27017b42,
        64'h7ae26a06_69a66946,
        64'h64e670a6_740600ff,
        64'hf797870e_c3c4c607,
        64'h87932481_00fff797,
        64'hc727a423_00fff797,
        64'h29010019_69138082,
        64'h6165853e_7b427ae2,
        64'h6a0669a6_694664e6,
        64'h740670a6_cd0187aa,
        64'h99028526_c9a58593,
        64'h009a1613_06a60dff,
        64'hf5974146_86b30019,
        64'h86934a01_05f00993,
        64'ha02169e2_6a4200fb,
        64'h08630081_6783fafb,
        64'h43e30b05_00816783,
        64'h08f70e63_770282e7,
        64'hb7830000_1797e531,
        64'h87aa9902_00faec63,
        64'h8f998a3a_89be0137,
        64'hf36305f7_0993000b,
        64'h186367e2_6742e7b5,
        64'h8526100c_862246c1,
        64'h87aa9902_02040613,
        64'h943e8526_080c0426,
        64'h036787b3_46c16402,
        64'h00c16783_05f00a93,
        64'h4b01cfad_4a0105f0,
        64'h099347a2_e14d87aa,
        64'h99028526_858a2480,
        64'h061346c1_08f71863,
        64'h89a7b783_77020000,
        64'h1797ed51_99028526,
        64'h100c2000_061346a1,
        64'h892af85a_fc56e0d2,
        64'he4cef0a2_f486e8ca,
        64'h84aeeca6_71598082,
        64'h4501b1ad_c291b37d,
        64'h4d81d71c_479ddfed,
        64'h01f7d79b_4b5cd35c,
        64'h000d3703_014d2783,
        64'hb54988d6_e002b3f9,
        64'h02100d93_bbd10200,
        64'h0d93bf59_6de2faeb,
        64'h05e32000_0713bf85,
        64'hf55fe0ef_417b0633,
        64'h65c2bfb5_f61fe0ef,
        64'h8556088c_865abbfd,
        64'hdc0d83e3_00050d9b,
        64'ha37ff0ef_f4bef882,
        64'hec82856a_08904785,
        64'h4685f0be_02610793,
        64'hc8be4791_e882b51d,
        64'h4de5b5d5_05010893,
        64'he03e4785_060b8563,
        64'h04940b63_bddd4d85,
        64'h05010893_e06eeeeb,
        64'h0fe32000_0713b5b9,
        64'h8daab55f_f0ef856a,
        64'h04c58593_46051034,
        64'h470115a2_06100593,
        64'h0af40263_4785ed84,
        64'h16e3200a_8a930c05,
        64'h060d9f63_bf91fc3e,
        64'he482e082_67a2d43e,
        64'h4789b569_4d81a821,
        64'hffdfe0ef_41760633,
        64'h20000613_65c20a0d,
        64'h9863015b_8533c795,
        64'h67820ce6_1d639341,
        64'h17420261_56038f55,
        64'h0086d69b_0086971b,
        64'hff9a10e3_8eb90c85,
        64'h92c116c2_00075703,
        64'h972e837d_17028f31,
        64'h0086969b_0086d61b,
        64'h000cc703_e4c18593,
        64'h4681ed49_2501b1df,
        64'hf0efe0ba_e482f802,
        64'h856a1030_47094685,
        64'hfc3a0261_0713d43a,
        64'h010d2583_4711f402,
        64'hfd3a1de3_e1711009,
        64'h89932501_b4bff0ef,
        64'h856a1030_4685010d,
        64'h2583e0a6_fc4ed44a,
        64'he4820a09_8663f802,
        64'hf4021000_04934911,
        64'h89c62008_8a138cc6,
        64'he00288d6_10ec0163,
        64'hfff40713_100c0e63,
        64'h18e69163_0fe00713,
        64'hb785fc0d_8ae33cfd,
        64'h00050d9b_b9bff0ef,
        64'he0a6fc4a_d44ee482,
        64'hf802856a_10304685,
        64'hf402010d_25830346,
        64'h95630251_4683160c,
        64'h8463a039_0ff00a13,
        64'h44850251_09134991,
        64'h71070c93_6709e83e,
        64'h4c01417a_8ab397de,
        64'h089ce43e_800c8793,
        64'hec3e6c85_017037b3,
        64'hb5fd0510_05938082,
        64'h2c010113_25813d83,
        64'h856e2601_3d032681,
        64'h3c832701_3c032781,
        64'h3b832801_3b032881,
        64'h3a832901_3a032981,
        64'h39832a01_39032a81,
        64'h34832b01_34032b81,
        64'h30834dc9_f8f1000d,
        64'h946334fd_00050d9b,
        64'hc3fff0ef_f4caf0ce,
        64'hc8d2f882_ec82856a,
        64'h08904685_e882010d,
        64'h25830607_d7630251,
        64'h0783a029_49050251,
        64'h09934a11_44a120f7,
        64'h0e63010d_258304c0,
        64'h07930281_4703040d,
        64'h98630005_0d9bc85f,
        64'hf0eff4be_f882ec82,
        64'h856a0890_47994685,
        64'hf0be103c_c8be478d,
        64'h010d2583_f43ee882,
        64'h8fd117a2_0017e793,
        64'h00171793_fed515e3,
        64'h0007c703_97ae0ff7,
        64'hf7938fb9_06850017,
        64'h171b0006_c78304c1,
        64'h85934701_05510513,
        64'h0894e8b2_8e4d8e5d,
        64'h8ff99381_076257fd,
        64'h8e5d8e75_0086571b,
        64'h00ff06b7_8fd507a2,
        64'h16820ff6_76930186,
        64'h579b8225_05200593,
        64'h10f40b63_47852404,
        64'h0a6302f1_02a38025,
        64'hfaa00793_945e1ff6,
        64'h84132000_0b13000b,
        64'h14631ff6_7b938aae,
        64'h8d2a1ffb_7b1325b1,
        64'h3c232791_34232781,
        64'h38232941_38232931,
        64'h3c232b21_30232a91,
        64'h34232a81_38232a11,
        64'h3c2327a1_30232771,
        64'h3c232951_342300d6,
        64'h0b332961_3023d401,
        64'h01138082_61450007,
        64'h851b6942_64e28ff5,
        64'h740270a2_80826145,
        64'h694264e2_740270a2,
        64'he7198f7d_0126c733,
        64'h37fd00e7_97bb0037,
        64'h171b4785_66a26398,
        64'h97b214c1_879301d7,
        64'h56130204_1713c485,
        64'he50de8df_f0ef8432,
        64'hf406f022_47010034,
        64'h893a84b6_e84aec26,
        64'h7179b725_444db735,
        64'h843edfe1_34fd0005,
        64'h079bde1f_f0eff852,
        64'hf456cc5a_fc02f002,
        64'h854e0830_4685ec02,
        64'h0109a583_f3c90171,
        64'h4783c49d_a0294a05,
        64'h01710a93_4b117104,
        64'h84936489_b7add81d,
        64'h0005041b_e1bff0ef,
        64'hf83efc02_f002854e,
        64'h08304785_4685f43e,
        64'h01710793_cc3e4791,
        64'hec02bf41_842ad171,
        64'h2501e41f_f0eff83e,
        64'hf452cc5e_fc02f002,
        64'h854e0830_46850a05,
        64'hec020109_a583bf55,
        64'h4401d71c_479ddfed,
        64'h01f7d79b_4b5cd35c,
        64'h0009b703_0149a783,
        64'hfc0918e3_e38517fd,
        64'h075b0863_639c97ba,
        64'h01d6d713_14c18793,
        64'h020b1693_80826149,
        64'h6ba66b46_6ae67a06,
        64'h79a67946_74e6640a,
        64'h852260aa_4449f8f9,
        64'he01934fd_0005041b,
        64'heb7ff0ef_f856f452,
        64'hcc5efc02_f002854e,
        64'h08304685_ec020109,
        64'ha5830407_d163000a,
        64'h0783a029_4a854b91,
        64'h44a10af7_06630109,
        64'ha58304c0_07930081,
        64'h4703e421_0005041b,
        64'hef7ff0ef_f83efc02,
        64'hf002893a_89aae4de,
        64'hecd6fca6_e506f4ce,
        64'hf8cae122_46850830,
        64'h8a364799_8b32f43e,
        64'he8daf0d2_003ccc3e,
        64'h490c478d_ec02e42e,
        64'h7175bfb9_d71c2781,
        64'h2007e793_8fd58ef1,
        64'h1ff7f793_c0060613,
        64'h00a6969b_37fd6605,
        64'h44140104_5783bf79,
        64'h450db759_d71c2007,
        64'h87936789_609802f7,
        64'h08230084_4783fed7,
        64'h8de30ff7_f7934b5c,
        64'h04800693_80826105,
        64'h450164a2_644260e2,
        64'hc01ff0ef_8526680c,
        64'h01845603_fce795e3,
        64'h4711401c_f1752501,
        64'hb75ff0ef_852685a2,
        64'h460104f6_ea6337f5,
        64'h80826105_64a26442,
        64'h60e24501_c35ff0ef,
        64'h85266c0c_02045603,
        64'h04e79263_471502e7,
        64'h8f634711_401ca93f,
        64'hf0ef8526_85a24601,
        64'hc3bd02f6_eb6308d7,
        64'h8a634689_401cdfed,
        64'h01f7d79b_4b5cd34c,
        64'h843284aa_ec06e426,
        64'he8221101_6118bf4d,
        64'h4555b5ed_470dd808,
        64'hbf41d41c_27818fd9,
        64'h1ff77713_8fd1377d,
        64'h0096161b_8ff500a7,
        64'h979b40c9_863b66c2,
        64'h010a5703_008a2783,
        64'h80826115_7dea6d0e,
        64'h6cae6c4e_6bee7b0e,
        64'h7aae7a4e_79ee6912,
        64'h64b26452_60f2450d,
        64'ha0112501_dd712501,
        64'hc35ff0ef_856a85d2,
        64'h00ebea63_3775b739,
        64'h000a2703_000d3403,
        64'hf96a82e3_028a0a13,
        64'h0a85d71c_27810127,
        64'he7b3000d_370302e4,
        64'h08230097_979b40c9,
        64'h87bb008a_4703ff97,
        64'h8de30ff7_f793485c,
        64'ha8914501_eefc63e3,
        64'h100c0c13_67a2ffbc,
        64'h93e3d33f_f0ef028d,
        64'h8d93856a_010db583,
        64'h018dd603_ff2791e3,
        64'h000da783_03bc8163,
        64'h028d8d93_d55ff0ef,
        64'h018db583_020dd603,
        64'h00879863_856aa831,
        64'h44154911_078d8c93,
        64'h096a9263_028a0a13,
        64'h0a85d41c_27810127,
        64'he7b38fd9_8fd18ff5,
        64'h0096161b_00a7979b,
        64'h40c9863b_66c2008a,
        64'h27834709_d8080085,
        64'h551b1097_8f636662,
        64'h00ca2783_e48ff0ef,
        64'hec32010a_2503ff97,
        64'h8de30ff7_f793485c,
        64'hc34d0eeb_e0631177,
        64'h0d63dfed_01f7d79b,
        64'h485c0016_3613ffea,
        64'h86134b0d_69090480,
        64'h0c934b89_4a814701,
        64'h8a6ed058_f13e0381,
        64'h0d93000d_3403010d,
        64'h27031000_079300f7,
        64'h74631000_07134187,
        64'h87b3d6a6_d0a604d1,
        64'h0023f502_e902e102,
        64'hfc82ec82_e882e482,
        64'hfc02c53a_4711d8ba,
        64'h46cde502_67a2ed3e,
        64'h97e2f482_f0827782,
        64'h00fc073b_e082f882,
        64'h77a24985_e83e4485,
        64'h8d2ac00a_87936a85,
        64'h12078863_4c0167a2,
        64'h1ce7ed63_e436f432,
        64'hf02e07f7_8793fd6e,
        64'he1eae5e6_e9e2edde,
        64'hf1daf5d6_f9d2fdce,
        64'he24ae626_ea22ee06,
        64'h02faf7b7_712d6518,
        64'hbddd86ae_8082450d,
        64'hbf01268d_feb81be3,
        64'h0087d79b_058500f5,
        64'h84239836_00d105b3,
        64'h00410813_80824501,
        64'he20dbf0d_268d4682,
        64'hfef6ac23_968a06c1,
        64'he9992781_0036f593,
        64'h55dcdbfd_0ff7f793,
        64'h0087d79b_49dc610c,
        64'hbf0dfe68_1be30087,
        64'hd79b0805_00f80423,
        64'h933a00e1_08330041,
        64'h0313b7b1_4702fef7,
        64'h2c23970a_07410008,
        64'h18632781_00377813,
        64'h02c82783_dbf50ff7,
        64'hf7930087_d79b0148,
        64'h27830005_3803bf2d,
        64'h270dff06_9be30087,
        64'hd79b0685_00f68423,
        64'h983a00e1_06b30041,
        64'h0813bf99_270d4702,
        64'hfef72c23_970a0741,
        64'hea812781_00377693,
        64'h56dcdbfd_0ff7f793,
        64'h0087d79b_4adc6114,
        64'h80820141_4501fef6,
        64'h11e393c1_03071793,
        64'he43e83a1_67a2fef7,
        64'h0fa3c036_07050081,
        64'h478336fd_0ad05863,
        64'h92411642_46829e39,
        64'h8736c61d_8a0dfed5,
        64'h96e30591_c43e0105,
        64'ha023c03a_47b24822,
        64'h377108e8_d863488d,
        64'h96be0045_8793068a,
        64'h470292c9_16c2ffc6,
        64'h069b12c7_fd63478d,
        64'hfff19241_0035f793,
        64'he43e83a1_c03a1642,
        64'h67a2fef5_8fa3367d,
        64'h05850081_4783377d,
        64'h08e05663_c6414701,
        64'hc78d0035_f793e402,
        64'he0021141_14058763,
        64'h16050a63_bf79678d,
        64'hebdff0ef_86260087,
        64'ha903698c_0205d483,
        64'hbf4d6789_ed1ff0ef,
        64'h86260087_a903698c,
        64'h0185d483_80826145,
        64'h450169a2_694264e2,
        64'hd71c2781_8fc57402,
        64'h70a21ff4_f4930127,
        64'he7b30009_b70334fd,
        64'h8fc100e9_793300a9,
        64'h191bc007_07130094,
        64'h141b6705_00144413,
        64'h67850185_d4830085,
        64'ha9038082_6145450d,
        64'h69a26942_64e27402,
        64'h70a204d7_0d63468d,
        64'h06d70a63_469502d7,
        64'h00638432_89aa87ae,
        64'h4691e84a_ec26f406,
        64'he44ef022_71794198,
        64'h80824501_fef712e3,
        64'h03068823_93c10305,
        64'h97930585_0005c803,
        64'hfec78de3_0ff7f793,
        64'h4adc6114_93410480,
        64'h06131742_00c8073b,
        64'hde5d85c2_8a0dff05,
        64'h98e3db1c_0591419c,
        64'hfed78de3_0ff7f793,
        64'h4b5c0480_0693983e,
        64'h00458793_080a6118,
        64'h03285813_1842ffc6,
        64'h081b02c7_f963882e,
        64'h478d8082_450dde75,
        64'h80824501_fe79c799,
        64'h92410035_f7931642,
        64'h02f70823_0585367d,
        64'h0005c783_fed78de3,
        64'h0ff7f793_4b5c6118,
        64'hc21d0480_0693cb9d,
        64'h0035f793_c99dcd0d,
        64'hb7e9468d_d8088082,
        64'h61056902_64a26442,
        64'hd41c60e2_27818fd9,
        64'h67098fd9_0096e733,
        64'h8ff900a7_979bc007,
        64'h07130094_949b6705,
        64'h0014c493_00892783,
        64'h4689d808_0085551b,
        64'h02f70f63_478500c9,
        64'h2703a37f_f0ef0109,
        64'h2503fee7_8de30ff7,
        64'hf793485c_04800713,
        64'h84b2892e_ec06e04a,
        64'he4266100_e8221101,
        64'h80820005_2823fbf5,
        64'h0ff7f793_8fd90087,
        64'hd71b495c_ffe58b85,
        64'h01e7d79b_495cc91c,
        64'h400007b7_bd554522,
        64'hfec710e3_070590d7,
        64'h87230100_2797dbe5,
        64'h0207f793_0147c783,
        64'h92078793_01002797,
        64'h00074683_00380070,
        64'h92e78823_01002797,
        64'h4751dbe5_0207f793,
        64'h0147c783_94478793,
        64'h01002797_0ff0000f,
        64'hc42a9782_0000100f,
        64'h67820ff0_000f96e7,
        64'h80234719_01002797,
        64'hdbe50207_f7930147,
        64'hc7839727_87930100,
        64'h2797ea1f_f0ef850a,
        64'h45a1b711_98878223,
        64'h01002797_dbe50207,
        64'hf7930147_c7839967,
        64'h87930100_2797fee6,
        64'h10e30705_9ad78223,
        64'h01002797_dbe50207,
        64'hf7930147_c7839b67,
        64'h87930100_27970007,
        64'h4683963a_c6056702,
        64'h9c978423_01002797,
        64'h6622dbe5_0207f793,
        64'h0147c783_9dc78793,
        64'h01002797_f0bff0ef,
        64'h002845a1_f13ff0ef,
        64'h850a45a1_bf9d9e87,
        64'h8b230100_2797dbe5,
        64'h0207f793_0147c783,
        64'ha0878793_01002797,
        64'hf37ff0ef_a0978a23,
        64'h01002797_650265a2,
        64'hdbe50207_f7930147,
        64'hc783a2a7_87930100,
        64'h2797f59f_f0ef0028,
        64'h45a1f61f_f0ef850a,
        64'h45a18082_61216a42,
        64'h69e27902_74a27442,
        64'h70e24505_07278263,
        64'h0d378d63_01470f63,
        64'h0ff77793_a647c703,
        64'h01002797_dbed8b85,
        64'h0147c783_a7478793,
        64'h01002797_0ff0000f,
        64'h494549cd_44114499,
        64'h4a49a8e7_86234719,
        64'h01002797_dbe50207,
        64'hf7930147_c783a9e7,
        64'h87930100_2797e852,
        64'hec4ef04a_f426f822,
        64'hfc067139_8082fee5,
        64'h11e3fef5_0fa30505,
        64'hac07c783_01002797,
        64'hdbed8b85_0147c783,
        64'had078793_01002797,
        64'h00b50733_c5858082,
        64'h0141450d_a011c31c,
        64'h00d80733_27819281,
        64'h8fd91682_8fd10187,
        64'h171b8b3d_0146161b,
        64'h0008b803_8fcd0108,
        64'h159b8a3d_8fcd0067,
        64'he7b300f8_781301f3,
        64'h131b01c7_e7b300a1,
        64'h470301de_1e1b01e7,
        64'h979b0091_46030081,
        64'h480300d1_430300b1,
        64'h4e0300c1_4783ed31,
        64'h0007851b_8fed35fd,
        64'h0015d59b_0026969b,
        64'h269988aa_77c102f5,
        64'hd5bbcfa5_4782cdb5,
        64'h9581c141_e432e02e,
        64'h1141bfe1_d54ddb5f,
        64'hf0ef86a2_47014087,
        64'h84330400_0793b7f5,
        64'h45018082_61216aa2,
        64'h6a4269e2_790274a2,
        64'h744270e2_dd71dddf,
        64'hf0ef0400_069300da,
        64'hf4630404_0413854e,
        64'h4701008a_05b30089,
        64'h06334084_86b30294,
        64'h7c63a82d_00946563,
        64'h04000a93_e42184b6,
        64'h8a2e89aa_893203f6,
        64'h7413e456_fc06e852,
        64'hec4ef04a_f426f822,
        64'h7139bd99_19019aca,
        64'h99caf52c_7ce3c89c,
        64'h0017e793_1b81489c,
        64'hffb90005_079bde5f,
        64'hf0ef8522_46054685,
        64'h0007c583_017987b3,
        64'hbfb5ff39_18e30985,
        64'h00f98023_00098463,
        64'h27814f9c_601c994e,
        64'hff27ebe3_07f7f793,
        64'h0107d79b_50dcc89c,
        64'h0017e793_489cf3d5,
        64'h0005079b_e2bff0ef,
        64'h85220ff9_7593460d,
        64'h4681ffc5_0005079b,
        64'he3fff0ef_85220a10,
        64'h05934601_4685f7f1,
        64'h0005079b_e53ff0ef,
        64'h85224609_46858082,
        64'h61656ce2_85666da2,
        64'h6d427c02_7ba27b42,
        64'h7ae26a06_69a66946,
        64'h64e67406_70a64c8d,
        64'ha0118cbe_d3f50d85,
        64'h0005079b_e8bff0ef,
        64'h85224605_46850007,
        64'hc58301b9_87b30bad,
        64'hf563a075_000b9563,
        64'h4d810200_0d13017c,
        64'h74638d5e_eb8d0005,
        64'h079beb9f_f0ef8522,
        64'h46054685_060b0563,
        64'h0ffaf593_040c9963,
        64'h00050c9b_ed3ff0ef,
        64'h85220ff5_f5934605,
        64'h4685008a_d593060c,
        64'h96630005_0c9beedf,
        64'hf0ef8522_0a000593,
        64'hc89c9bf9_46014685,
        64'h489cfcd7_eee38fd9,
        64'h93011702_1782ff85,
        64'h2703ffc7_a7839552,
        64'h97d2d365_0513d3a7,
        64'h87930004_05170004,
        64'h07970685_8edd9381,
        64'h17821682_ff87a783,
        64'hffc72683_97d29752,
        64'hd5c78793_d6070713,
        64'h00040797_00040717,
        64'hfff107f7_f7938fc9,
        64'h0187d79b_8d590087,
        64'hd51b0107_d71bf96d,
        64'h278107f7_f51350dc,
        64'h60040e04_0b630200,
        64'h0c136a31_fff68b93,
        64'h8b3a8ab2_89ae842a,
        64'h8936e46e_e86aec66,
        64'heca6f486_f062f45e,
        64'hf85afc56_e0d2e4ce,
        64'he8caf0a2_7159bf75,
        64'h46014705_4801b7d1,
        64'h47014805_4601fef5,
        64'h8082450d_faf76fe3,
        64'h4709ffd6_079b8082,
        64'h4501cedc_27818fd9,
        64'h0097171b_0107e7b3,
        64'h611400a8_181b8fd1,
        64'h0086161b_00d5e7b3,
        64'h00c6969b_47014801,
        64'h00c03633_167d04f6,
        64'h0163478d_04f60963,
        64'h4789ee9d_c5298082,
        64'hfca7eee3_8fd99301,
        64'h17021782_ff872703,
        64'hffc7a783_973697b6,
        64'he3c70713_e4078793,
        64'h00040717_00040797,
        64'h66b18082_fa6d0585,
        64'h0305167d_00730023,
        64'h00058383_ca09832a,
        64'h80822501_8d5d8d79,
        64'h00ff0737_0085151b,
        64'h8fd98f75_0085571b,
        64'hf0068693_8fd966c1,
        64'h0185579b_0185171b,
        64'hbff51050_007300a2,
        64'ha423e922_82930100,
        64'h02970015_65130506,
        64'h342010ef_0000100f,
        64'h0ff0000f_43014281,
        64'h80820002_80e7f140,
        64'h25730062_e2b30102,
        64'he2831302_0142e303,
        64'hec828293_01000297,
        64'hfe72cbe3_0291fe03,
        64'h1ee30002_a3039396,
        64'h038a04c3_a383ee63,
        64'h83930100_03970003,
        64'h20239316_030af140,
        64'h2373efa2_82930004,
        64'h0297fe03_0ae30083,
        64'h73133440_23731050,
        64'h0073fe72_cce30291,
        64'h0062a023_43059396,
        64'h038a04c3_a383f263,
        64'h83930100_0397f2e2,
        64'h82930004_02970ff0,
        64'h000f00a2_aa239101,
        64'h00a2a823_f4428293,
        64'h01000297_92820a02,
        64'h81630482_a283f562,
        64'h82930100_02971161,
        64'h91160542_a283f661,
        64'h01130e00_0117f6e2,
        64'h82930100_02970062,
        64'ha8234305_0062a223,
        64'h0062a023_537dfe03,
        64'h0ee30482_a303f8e2,
        64'h82930100_12970202,
        64'h8e630022_f2930502,
        64'ha283fa22_82930100,
        64'h029798e1_81930000,
        64'h2197faa1_01130e01,
        64'h01170a62_9663f140,
        64'h23734281_30431073,
        64'h43214f81_4f014e81,
        64'h4e014d81_4d014c81,
        64'h4c014b81_4b014a81,
        64'h4a014981_49014881,
        64'h48014781_47014681,
        64'h46014581_45014481,
        64'h44014381_43014281,
        64'h42014181_41014081
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
