// Copyright 2020 ETH Zurich
    // SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
    //
    // Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
    // Florian Zaruba <zarubaf@iis.ee.ethz.ch>
    // Stefan Mach <smach@iis.ee.ethz.ch>
    // Thomas Benz <tbenz@iis.ee.ethz.ch>
    // Paul Scheffler <paulsc@iis.ee.ethz.ch>
    // Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
    //
    // AUTOMATICALLY GENERATED by gen_bootrom.py; edit the script instead.

    module bootrom #(
        parameter int unsigned AddrWidth = 32,
        parameter int unsigned DataWidth = 32
    )(
        input  logic                 clk_i,
        input  logic                 rst_ni,
        input  logic                 req_i,
        input  logic [AddrWidth-1:0] addr_i,
        output logic [DataWidth-1:0] data_o
    );
        localparam NumWords   = 16384;
        logic [$clog2(NumWords)-1:0] word;

        assign word = addr_i / (DataWidth / 8);

        always_comb begin
            data_o = '0;
            unique case (word)
                000: data_o = 32'h6f020117 /* 0x0000 */;
                001: data_o = 32'hff810113 /* 0x0004 */;
                002: data_o = 32'h00000197 /* 0x0008 */;
                003: data_o = 32'h59918193 /* 0x000c */;
                004: data_o = 32'h42014081 /* 0x0010 */;
                005: data_o = 32'h43014281 /* 0x0014 */;
                006: data_o = 32'h44014381 /* 0x0018 */;
                007: data_o = 32'h45014481 /* 0x001c */;
                008: data_o = 32'h46014581 /* 0x0020 */;
                009: data_o = 32'h47014681 /* 0x0024 */;
                010: data_o = 32'h48014781 /* 0x0028 */;
                011: data_o = 32'h49014881 /* 0x002c */;
                012: data_o = 32'h4a014981 /* 0x0030 */;
                013: data_o = 32'h4b014a81 /* 0x0034 */;
                014: data_o = 32'h4c014b81 /* 0x0038 */;
                015: data_o = 32'h4d014c81 /* 0x003c */;
                016: data_o = 32'h4e014d81 /* 0x0040 */;
                017: data_o = 32'h4f014e81 /* 0x0044 */;
                018: data_o = 32'h0000100f /* 0x0048 */;
                019: data_o = 32'h280000ef /* 0x004c */;
                020: data_o = 32'h0506a009 /* 0x0050 */;
                021: data_o = 32'h00156513 /* 0x0054 */;
                022: data_o = 32'h020042b7 /* 0x0058 */;
                023: data_o = 32'h00a2a223 /* 0x005c */;
                024: data_o = 32'h10500073 /* 0x0060 */;
                025: data_o = 32'h0617bff5 /* 0x0064 */;
                026: data_o = 32'h71190200 /* 0x0068 */;
                027: data_o = 32'hf9a60613 /* 0x006c */;
                028: data_o = 32'hf8a6fca2 /* 0x0070 */;
                029: data_o = 32'hf0cef4ca /* 0x0074 */;
                030: data_o = 32'he8d6ecd2 /* 0x0078 */;
                031: data_o = 32'h87aae4da /* 0x007c */;
                032: data_o = 32'h86b24741 /* 0x0080 */;
                033: data_o = 32'he58396ba /* 0x0084 */;
                034: data_o = 32'hde2e0006 /* 0x0088 */;
                035: data_o = 32'h053756f2 /* 0x008c */;
                036: data_o = 32'h85b28000 /* 0x0090 */;
                037: data_o = 32'hdc362681 /* 0x0094 */;
                038: data_o = 32'h8ec956e2 /* 0x0098 */;
                039: data_o = 32'h56e2dc36 /* 0x009c */;
                040: data_o = 32'hc19495ba /* 0x00a0 */;
                041: data_o = 32'h000c36b7 /* 0x00a4 */;
                042: data_o = 32'h50068693 /* 0x00a8 */;
                043: data_o = 32'h02d7d7b3 /* 0x00ac */;
                044: data_o = 32'h0fff05b7 /* 0x00b0 */;
                045: data_o = 32'h37fd86b2 /* 0x00b4 */;
                046: data_o = 32'h0107979b /* 0x00b8 */;
                047: data_o = 32'h0107d79b /* 0x00bc */;
                048: data_o = 32'h45e18fcd /* 0x00c0 */;
                049: data_o = 32'hc29c96ae /* 0x00c4 */;
                050: data_o = 32'h87b24681 /* 0x00c8 */;
                051: data_o = 32'h02000593 /* 0x00cc */;
                052: data_o = 32'hc39497ae /* 0x00d0 */;
                053: data_o = 32'h97ba87b2 /* 0x00d4 */;
                054: data_o = 32'h0007e683 /* 0x00d8 */;
                055: data_o = 32'h57d2da36 /* 0x00dc */;
                056: data_o = 32'h278186b2 /* 0x00e0 */;
                057: data_o = 32'h57c2d83e /* 0x00e4 */;
                058: data_o = 32'hf7932781 /* 0x00e8 */;
                059: data_o = 32'he793f007 /* 0x00ec */;
                060: data_o = 32'hd83e0087 /* 0x00f0 */;
                061: data_o = 32'h96ba57c2 /* 0x00f4 */;
                062: data_o = 32'h0813c29c /* 0x00f8 */;
                063: data_o = 32'h00337d00 /* 0x00fc */;
                064: data_o = 32'h387d0000 /* 0x0100 */;
                065: data_o = 32'hfe081de3 /* 0x0104 */;
                066: data_o = 32'h6f000497 /* 0x0108 */;
                067: data_o = 32'h6909678d /* 0x010c */;
                068: data_o = 32'h6f000597 /* 0x0110 */;
                069: data_o = 32'hef848493 /* 0x0114 */;
                070: data_o = 32'h02000517 /* 0x0118 */;
                071: data_o = 32'h10078793 /* 0x011c */;
                072: data_o = 32'h0a9b6985 /* 0x0120 */;
                073: data_o = 32'h85932009 /* 0x0124 */;
                074: data_o = 32'h94beff05 /* 0x0128 */;
                075: data_o = 32'hf1050513 /* 0x012c */;
                076: data_o = 32'h04134751 /* 0x0130 */;
                077: data_o = 32'h091b0240 /* 0x0134 */;
                078: data_o = 32'h899b2029 /* 0x0138 */;
                079: data_o = 32'h6a410ff9 /* 0x013c */;
                080: data_o = 32'h00386793 /* 0x0140 */;
                081: data_o = 32'h87b2c11c /* 0x0144 */;
                082: data_o = 32'he68397ba /* 0x0148 */;
                083: data_o = 32'hc8360007 /* 0x014c */;
                084: data_o = 32'h278147c2 /* 0x0150 */;
                085: data_o = 32'h47b2c63e /* 0x0154 */;
                086: data_o = 32'h01f7d79b /* 0x0158 */;
                087: data_o = 32'h87b2d7ed /* 0x015c */;
                088: data_o = 32'ha02397a2 /* 0x0160 */;
                089: data_o = 32'h87b20157 /* 0x0164 */;
                090: data_o = 32'he68397ba /* 0x0168 */;
                091: data_o = 32'hcc360007 /* 0x016c */;
                092: data_o = 32'h278147e2 /* 0x0170 */;
                093: data_o = 32'h47d2ca3e /* 0x0174 */;
                094: data_o = 32'h01f7d79b /* 0x0178 */;
                095: data_o = 32'h87b2d7ed /* 0x017c */;
                096: data_o = 32'ha02397a2 /* 0x0180 */;
                097: data_o = 32'h87b20127 /* 0x0184 */;
                098: data_o = 32'he68397ba /* 0x0188 */;
                099: data_o = 32'hd0360007 /* 0x018c */;
                100: data_o = 32'h27815782 /* 0x0190 */;
                101: data_o = 32'h47f2ce3e /* 0x0194 */;
                102: data_o = 32'h01f7d79b /* 0x0198 */;
                103: data_o = 32'h87b2d7ed /* 0x019c */;
                104: data_o = 32'ha02397a2 /* 0x01a0 */;
                105: data_o = 32'h87b20137 /* 0x01a4 */;
                106: data_o = 32'he68397ba /* 0x01a8 */;
                107: data_o = 32'hd4360007 /* 0x01ac */;
                108: data_o = 32'h278157a2 /* 0x01b0 */;
                109: data_o = 32'h5792d23e /* 0x01b4 */;
                110: data_o = 32'h01f7d79b /* 0x01b8 */;
                111: data_o = 32'h8b13d7ed /* 0x01bc */;
                112: data_o = 32'h87b2f005 /* 0x01c0 */;
                113: data_o = 32'he68397ba /* 0x01c4 */;
                114: data_o = 32'hd6360007 /* 0x01c8 */;
                115: data_o = 32'h969357b2 /* 0x01cc */;
                116: data_o = 32'hd8e302b7 /* 0x01d0 */;
                117: data_o = 32'h6883fe06 /* 0x01d4 */;
                118: data_o = 32'h62830005 /* 0x01d8 */;
                119: data_o = 32'h63030005 /* 0x01dc */;
                120: data_o = 32'h63830005 /* 0x01e0 */;
                121: data_o = 32'h6e030005 /* 0x01e4 */;
                122: data_o = 32'h6e830005 /* 0x01e8 */;
                123: data_o = 32'h6f030005 /* 0x01ec */;
                124: data_o = 32'h6f830005 /* 0x01f0 */;
                125: data_o = 32'h20230005 /* 0x01f4 */;
                126: data_o = 32'h2223011b /* 0x01f8 */;
                127: data_o = 32'h2423005b /* 0x01fc */;
                128: data_o = 32'h2623006b /* 0x0200 */;
                129: data_o = 32'h2823007b /* 0x0204 */;
                130: data_o = 32'h2a2301cb /* 0x0208 */;
                131: data_o = 32'h2c2301db /* 0x020c */;
                132: data_o = 32'h2e2301eb /* 0x0210 */;
                133: data_o = 32'h0b1301fb /* 0x0214 */;
                134: data_o = 32'h94e3020b /* 0x0218 */;
                135: data_o = 32'h8593fb65 /* 0x021c */;
                136: data_o = 32'h083b1005 /* 0x0220 */;
                137: data_o = 32'h9de3010a /* 0x0224 */;
                138: data_o = 32'h100ff0b4 /* 0x0228 */;
                139: data_o = 32'h74660000 /* 0x022c */;
                140: data_o = 32'h792674c6 /* 0x0230 */;
                141: data_o = 32'h6a667986 /* 0x0234 */;
                142: data_o = 32'h6b266ac6 /* 0x0238 */;
                143: data_o = 32'h6f000597 /* 0x023c */;
                144: data_o = 32'hdc458593 /* 0x0240 */;
                145: data_o = 32'h61094501 /* 0x0244 */;
                146: data_o = 32'h6f000317 /* 0x0248 */;
                147: data_o = 32'hdb830067 /* 0x024c */;
                148: data_o = 32'hc691882a /* 0x0250 */;
                149: data_o = 32'hffd6079b /* 0x0254 */;
                150: data_o = 32'h75634509 /* 0x0258 */;
                151: data_o = 32'h479506f5 /* 0x025c */;
                152: data_o = 32'h04c7e863 /* 0x0260 */;
                153: data_o = 32'hfeb18793 /* 0x0264 */;
                154: data_o = 32'h963e060a /* 0x0268 */;
                155: data_o = 32'h97ba4218 /* 0x026c */;
                156: data_o = 32'h45098782 /* 0x0270 */;
                157: data_o = 32'h47858082 /* 0x0274 */;
                158: data_o = 32'h863efeed /* 0x0278 */;
                159: data_o = 32'h47814701 /* 0x027c */;
                160: data_o = 32'h969b4505 /* 0x0280 */;
                161: data_o = 32'h8dd500c6 /* 0x0284 */;
                162: data_o = 32'h36838dd9 /* 0x0288 */;
                163: data_o = 32'h979b0008 /* 0x028c */;
                164: data_o = 32'h8fcd0097 /* 0x0290 */;
                165: data_o = 32'h00a5151b /* 0x0294 */;
                166: data_o = 32'h161b8fc9 /* 0x0298 */;
                167: data_o = 32'h873600b6 /* 0x029c */;
                168: data_o = 32'h46f18fd1 /* 0x02a0 */;
                169: data_o = 32'hc31c9736 /* 0x02a4 */;
                170: data_o = 32'h80824501 /* 0x02a8 */;
                171: data_o = 32'hb7e94781 /* 0x02ac */;
                172: data_o = 32'h47054781 /* 0x02b0 */;
                173: data_o = 32'h0087171b /* 0x02b4 */;
                174: data_o = 32'h45014601 /* 0x02b8 */;
                175: data_o = 32'h4781b7d9 /* 0x02bc */;
                176: data_o = 32'hbfcd4701 /* 0x02c0 */;
                177: data_o = 32'h47858082 /* 0x02c4 */;
                178: data_o = 32'hb7ed4701 /* 0x02c8 */;
                179: data_o = 32'h01004797 /* 0x02cc */;
                180: data_o = 32'hd3478793 /* 0x02d0 */;
                181: data_o = 32'h711d4bdc /* 0x02d4 */;
                182: data_o = 32'he8a2ec86 /* 0x02d8 */;
                183: data_o = 32'he0cae4a6 /* 0x02dc */;
                184: data_o = 32'hf852fc4e /* 0x02e0 */;
                185: data_o = 32'h4709f456 /* 0x02e4 */;
                186: data_o = 32'h81632781 /* 0x02e8 */;
                187: data_o = 32'h6d630ee7 /* 0x02ec */;
                188: data_o = 32'h866300f7 /* 0x02f0 */;
                189: data_o = 32'hf5371007 /* 0x02f4 */;
                190: data_o = 32'h051302fa /* 0x02f8 */;
                191: data_o = 32'hf0ef0805 /* 0x02fc */;
                192: data_o = 32'h0073d69f /* 0x0300 */;
                193: data_o = 32'hbff51050 /* 0x0304 */;
                194: data_o = 32'h9c63470d /* 0x0308 */;
                195: data_o = 32'h27170ae7 /* 0x030c */;
                196: data_o = 32'h06b70100 /* 0x0310 */;
                197: data_o = 32'h07132201 /* 0x0314 */;
                198: data_o = 32'h8693cf27 /* 0x0318 */;
                199: data_o = 32'hc714d086 /* 0x031c */;
                200: data_o = 32'h01002717 /* 0x0320 */;
                201: data_o = 32'hc95806b7 /* 0x0324 */;
                202: data_o = 32'hce070713 /* 0x0328 */;
                203: data_o = 32'h19068693 /* 0x032c */;
                204: data_o = 32'h01001797 /* 0x0330 */;
                205: data_o = 32'h8793c354 /* 0x0334 */;
                206: data_o = 32'h0737cd07 /* 0x0338 */;
                207: data_o = 32'hec3e0104 /* 0x033c */;
                208: data_o = 32'h0787071b /* 0x0340 */;
                209: data_o = 32'h03000693 /* 0x0344 */;
                210: data_o = 32'hc39897b6 /* 0x0348 */;
                211: data_o = 32'h003c07b7 /* 0x034c */;
                212: data_o = 32'h879b66e2 /* 0x0350 */;
                213: data_o = 32'h06130c87 /* 0x0354 */;
                214: data_o = 32'h96b20340 /* 0x0358 */;
                215: data_o = 32'h07b7c29c /* 0x035c */;
                216: data_o = 32'h66e20078 /* 0x0360 */;
                217: data_o = 32'h0787879b /* 0x0364 */;
                218: data_o = 32'h03800613 /* 0x0368 */;
                219: data_o = 32'hc29c96b2 /* 0x036c */;
                220: data_o = 32'h66e267c1 /* 0x0370 */;
                221: data_o = 32'h061327d1 /* 0x0374 */;
                222: data_o = 32'h96b203c0 /* 0x0378 */;
                223: data_o = 32'h0693c29c /* 0x037c */;
                224: data_o = 32'h67e20400 /* 0x0380 */;
                225: data_o = 32'hc39897b6 /* 0x0384 */;
                226: data_o = 32'h67e24741 /* 0x0388 */;
                227: data_o = 32'he68397ba /* 0x038c */;
                228: data_o = 32'hc2360007 /* 0x0390 */;
                229: data_o = 32'h66e24792 /* 0x0394 */;
                230: data_o = 32'he7932781 /* 0x0398 */;
                231: data_o = 32'h96ba0017 /* 0x039c */;
                232: data_o = 32'h0824c29c /* 0x03a0 */;
                233: data_o = 32'h46014685 /* 0x03a4 */;
                234: data_o = 32'h0a000593 /* 0x03a8 */;
                235: data_o = 32'hf0ef8526 /* 0x03ac */;
                236: data_o = 32'h079bea3f /* 0x03b0 */;
                237: data_o = 32'hcbad0005 /* 0x03b4 */;
                238: data_o = 32'h10500073 /* 0x03b8 */;
                239: data_o = 32'h10500073 /* 0x03bc */;
                240: data_o = 32'h0073bfe5 /* 0x03c0 */;
                241: data_o = 32'h00731050 /* 0x03c4 */;
                242: data_o = 32'hbfe51050 /* 0x03c8 */;
                243: data_o = 32'h01002797 /* 0x03cc */;
                244: data_o = 32'h22010737 /* 0x03d0 */;
                245: data_o = 32'hc3478793 /* 0x03d4 */;
                246: data_o = 32'hd0870713 /* 0x03d8 */;
                247: data_o = 32'h2797c798 /* 0x03dc */;
                248: data_o = 32'h07370100 /* 0x03e0 */;
                249: data_o = 32'h8793c958 /* 0x03e4 */;
                250: data_o = 32'h0713c227 /* 0x03e8 */;
                251: data_o = 32'hc5371907 /* 0x03ec */;
                252: data_o = 32'h05130beb /* 0x03f0 */;
                253: data_o = 32'hc3d82005 /* 0x03f4 */;
                254: data_o = 32'hc6fff0ef /* 0x03f8 */;
                255: data_o = 32'h2797b719 /* 0x03fc */;
                256: data_o = 32'h07370100 /* 0x0400 */;
                257: data_o = 32'h87932201 /* 0x0404 */;
                258: data_o = 32'h0713c027 /* 0x0408 */;
                259: data_o = 32'hc798d087 /* 0x040c */;
                260: data_o = 32'h01002797 /* 0x0410 */;
                261: data_o = 32'hc9580737 /* 0x0414 */;
                262: data_o = 32'hbf078793 /* 0x0418 */;
                263: data_o = 32'h19070713 /* 0x041c */;
                264: data_o = 32'h0073c3d8 /* 0x0420 */;
                265: data_o = 32'hbff51050 /* 0x0424 */;
                266: data_o = 32'h46054685 /* 0x0428 */;
                267: data_o = 32'h85264581 /* 0x042c */;
                268: data_o = 32'he21ff0ef /* 0x0430 */;
                269: data_o = 32'h0005079b /* 0x0434 */;
                270: data_o = 32'h0073c781 /* 0x0438 */;
                271: data_o = 32'hbff51050 /* 0x043c */;
                272: data_o = 32'h46094685 /* 0x0440 */;
                273: data_o = 32'h85264581 /* 0x0444 */;
                274: data_o = 32'he09ff0ef /* 0x0448 */;
                275: data_o = 32'h0005079b /* 0x044c */;
                276: data_o = 32'h0073c781 /* 0x0450 */;
                277: data_o = 32'hbff51050 /* 0x0454 */;
                278: data_o = 32'h46014685 /* 0x0458 */;
                279: data_o = 32'h0a100593 /* 0x045c */;
                280: data_o = 32'hf0ef8526 /* 0x0460 */;
                281: data_o = 32'h079bdeff /* 0x0464 */;
                282: data_o = 32'heff10005 /* 0x0468 */;
                283: data_o = 32'h6f000417 /* 0x046c */;
                284: data_o = 32'h6f003917 /* 0x0470 */;
                285: data_o = 32'hb9440413 /* 0x0474 */;
                286: data_o = 32'hb5090913 /* 0x0478 */;
                287: data_o = 32'h02400a13 /* 0x047c */;
                288: data_o = 32'h03e00a93 /* 0x0480 */;
                289: data_o = 32'h468149e1 /* 0x0484 */;
                290: data_o = 32'h05934611 /* 0x0488 */;
                291: data_o = 32'h85260400 /* 0x048c */;
                292: data_o = 32'hdc1ff0ef /* 0x0490 */;
                293: data_o = 32'h0005079b /* 0x0494 */;
                294: data_o = 32'h67e2ebd5 /* 0x0498 */;
                295: data_o = 32'he70397d2 /* 0x049c */;
                296: data_o = 32'hc43a0007 /* 0x04a0 */;
                297: data_o = 32'hd79b47a2 /* 0x04a4 */;
                298: data_o = 32'hf7930107 /* 0x04a8 */;
                299: data_o = 32'hf6e307f7 /* 0x04ac */;
                300: data_o = 32'h87a2fefa /* 0x04b0 */;
                301: data_o = 32'h04040693 /* 0x04b4 */;
                302: data_o = 32'h974e6762 /* 0x04b8 */;
                303: data_o = 32'h00076603 /* 0x04bc */;
                304: data_o = 32'h4732c632 /* 0x04c0 */;
                305: data_o = 32'hc3992701 /* 0x04c4 */;
                306: data_o = 32'h00e78023 /* 0x04c8 */;
                307: data_o = 32'h95e30785 /* 0x04cc */;
                308: data_o = 32'h0413fed7 /* 0x04d0 */;
                309: data_o = 32'h18e30404 /* 0x04d4 */;
                310: data_o = 32'h4681fb24 /* 0x04d8 */;
                311: data_o = 32'h05934615 /* 0x04dc */;
                312: data_o = 32'h08280400 /* 0x04e0 */;
                313: data_o = 32'hd6dff0ef /* 0x04e4 */;
                314: data_o = 32'h0005079b /* 0x04e8 */;
                315: data_o = 32'h0713e3bd /* 0x04ec */;
                316: data_o = 32'h06930240 /* 0x04f0 */;
                317: data_o = 32'h67e203e0 /* 0x04f4 */;
                318: data_o = 32'he60397ba /* 0x04f8 */;
                319: data_o = 32'hc8320007 /* 0x04fc */;
                320: data_o = 32'hd79b47c2 /* 0x0500 */;
                321: data_o = 32'hf7930107 /* 0x0504 */;
                322: data_o = 32'hf6e307f7 /* 0x0508 */;
                323: data_o = 32'h3797fef6 /* 0x050c */;
                324: data_o = 32'h87936f00 /* 0x0510 */;
                325: data_o = 32'h46e1af27 /* 0x0514 */;
                326: data_o = 32'h04056762 /* 0x0518 */;
                327: data_o = 32'h66039736 /* 0x051c */;
                328: data_o = 32'hca320007 /* 0x0520 */;
                329: data_o = 32'h0fa34752 /* 0x0524 */;
                330: data_o = 32'h17e3fee4 /* 0x0528 */;
                331: data_o = 32'h100ffef4 /* 0x052c */;
                332: data_o = 32'h05970000 /* 0x0530 */;
                333: data_o = 32'h85936f00 /* 0x0534 */;
                334: data_o = 32'h4501ace5 /* 0x0538 */;
                335: data_o = 32'h6f000097 /* 0x053c */;
                336: data_o = 32'hac4080e7 /* 0x0540 */;
                337: data_o = 32'h0073bb7d /* 0x0544 */;
                338: data_o = 32'hbff51050 /* 0x0548 */;
                339: data_o = 32'h10500073 /* 0x054c */;
                340: data_o = 32'h0073bff5 /* 0x0550 */;
                341: data_o = 32'hbff51050 /* 0x0554 */;
                342: data_o = 32'h00003241 /* 0x0558 */;
                343: data_o = 32'h73697200 /* 0x055c */;
                344: data_o = 32'h01007663 /* 0x0560 */;
                345: data_o = 32'h00000028 /* 0x0564 */;
                346: data_o = 32'h36767205 /* 0x0568 */;
                347: data_o = 32'h70326934 /* 0x056c */;
                348: data_o = 32'h326d5f30 /* 0x0570 */;
                349: data_o = 32'h615f3070 /* 0x0574 */;
                350: data_o = 32'h5f307032 /* 0x0578 */;
                351: data_o = 32'h30703266 /* 0x057c */;
                352: data_o = 32'h7032645f /* 0x0580 */;
                353: data_o = 32'h32635f30 /* 0x0584 */;
                354: data_o = 32'h00003070 /* 0x0588 */;
                355: data_o = 32'hfffffd24 /* 0x058c */;
                356: data_o = 32'hfffffd32 /* 0x0590 */;
                357: data_o = 32'hfffffd3a /* 0x0594 */;
                358: data_o = 32'hfffffd20 /* 0x0598 */;
                359: data_o = 32'hfffffcea /* 0x059c */;
                360: data_o = 32'hfffffce6 /* 0x05a0 */;
                361: data_o = 32'h3a434347 /* 0x05a4 */;
                362: data_o = 32'h4e472820 /* 0x05a8 */;
                363: data_o = 32'h39202955 /* 0x05ac */;
                364: data_o = 32'h302e322e /* 0x05b0 */;
                365: data_o = 32'h00344100 /* 0x05b4 */;
                366: data_o = 32'h69720000 /* 0x05b8 */;
                367: data_o = 32'h00766373 /* 0x05bc */;
                368: data_o = 32'h00002a01 /* 0x05c0 */;
                369: data_o = 32'h05100400 /* 0x05c4 */;
                370: data_o = 32'h34367672 /* 0x05c8 */;
                371: data_o = 32'h30703269 /* 0x05cc */;
                372: data_o = 32'h70326d5f /* 0x05d0 */;
                373: data_o = 32'h32615f30 /* 0x05d4 */;
                374: data_o = 32'h665f3070 /* 0x05d8 */;
                375: data_o = 32'h5f307032 /* 0x05dc */;
                376: data_o = 32'h30703264 /* 0x05e0 */;
                377: data_o = 32'h7032635f /* 0x05e4 */;
                378: data_o = 32'h00000030 /* 0x05e8 */;
                379: data_o = 32'h00000000 /* 0x05ec */;
                380: data_o = 32'h00000000 /* 0x05f0 */;
                381: data_o = 32'h00000000 /* 0x05f4 */;
                382: data_o = 32'h00000000 /* 0x05f8 */;
                383: data_o = 32'h00000000 /* 0x05fc */;
                384: data_o = 32'h00000000 /* 0x0600 */;
                385: data_o = 32'h00000000 /* 0x0604 */;
                386: data_o = 32'h00000000 /* 0x0608 */;
                387: data_o = 32'h00000000 /* 0x060c */;
                388: data_o = 32'h00000000 /* 0x0610 */;
                389: data_o = 32'h00000000 /* 0x0614 */;
                390: data_o = 32'h00000000 /* 0x0618 */;
                391: data_o = 32'h00000000 /* 0x061c */;
                392: data_o = 32'h00000000 /* 0x0620 */;
                393: data_o = 32'h00000000 /* 0x0624 */;
                394: data_o = 32'h00000000 /* 0x0628 */;
                395: data_o = 32'h00000000 /* 0x062c */;
                396: data_o = 32'h00000000 /* 0x0630 */;
                397: data_o = 32'h00000000 /* 0x0634 */;
                398: data_o = 32'h00000000 /* 0x0638 */;
                399: data_o = 32'h00000000 /* 0x063c */;
                400: data_o = 32'h00000000 /* 0x0640 */;
                401: data_o = 32'h00000000 /* 0x0644 */;
                402: data_o = 32'h00000000 /* 0x0648 */;
                403: data_o = 32'h00000000 /* 0x064c */;
                404: data_o = 32'h00000000 /* 0x0650 */;
                405: data_o = 32'h00000000 /* 0x0654 */;
                406: data_o = 32'h00000000 /* 0x0658 */;
                407: data_o = 32'h00000000 /* 0x065c */;
                408: data_o = 32'h00000000 /* 0x0660 */;
                409: data_o = 32'h00000000 /* 0x0664 */;
                410: data_o = 32'h00000000 /* 0x0668 */;
                411: data_o = 32'h00000000 /* 0x066c */;
                412: data_o = 32'h00000000 /* 0x0670 */;
                413: data_o = 32'h00000000 /* 0x0674 */;
                414: data_o = 32'h00000000 /* 0x0678 */;
                415: data_o = 32'h00000000 /* 0x067c */;
                416: data_o = 32'h00000000 /* 0x0680 */;
                417: data_o = 32'h00000000 /* 0x0684 */;
                418: data_o = 32'h00000000 /* 0x0688 */;
                419: data_o = 32'h00000000 /* 0x068c */;
                420: data_o = 32'h00000000 /* 0x0690 */;
                421: data_o = 32'h00000000 /* 0x0694 */;
                422: data_o = 32'h00000000 /* 0x0698 */;
                423: data_o = 32'h00000000 /* 0x069c */;
                424: data_o = 32'h00000000 /* 0x06a0 */;
                425: data_o = 32'h00000000 /* 0x06a4 */;
                426: data_o = 32'h00000000 /* 0x06a8 */;
                427: data_o = 32'h00000000 /* 0x06ac */;
                428: data_o = 32'h00000000 /* 0x06b0 */;
                429: data_o = 32'h00000000 /* 0x06b4 */;
                430: data_o = 32'h00000000 /* 0x06b8 */;
                431: data_o = 32'h00000000 /* 0x06bc */;
                432: data_o = 32'h00000000 /* 0x06c0 */;
                433: data_o = 32'h00000000 /* 0x06c4 */;
                434: data_o = 32'h00000000 /* 0x06c8 */;
                435: data_o = 32'h00000000 /* 0x06cc */;
                436: data_o = 32'h00000000 /* 0x06d0 */;
                437: data_o = 32'h00000000 /* 0x06d4 */;
                438: data_o = 32'h00000000 /* 0x06d8 */;
                439: data_o = 32'h00000000 /* 0x06dc */;
                440: data_o = 32'h00000000 /* 0x06e0 */;
                441: data_o = 32'h00000000 /* 0x06e4 */;
                442: data_o = 32'h00000000 /* 0x06e8 */;
                443: data_o = 32'h00000000 /* 0x06ec */;
                444: data_o = 32'h00000000 /* 0x06f0 */;
                445: data_o = 32'h00000000 /* 0x06f4 */;
                446: data_o = 32'h00000000 /* 0x06f8 */;
                447: data_o = 32'h00000000 /* 0x06fc */;
                448: data_o = 32'h00000000 /* 0x0700 */;
                449: data_o = 32'h00000000 /* 0x0704 */;
                450: data_o = 32'h00000000 /* 0x0708 */;
                451: data_o = 32'h00000000 /* 0x070c */;
                452: data_o = 32'h00000000 /* 0x0710 */;
                453: data_o = 32'h00000000 /* 0x0714 */;
                454: data_o = 32'h00000000 /* 0x0718 */;
                455: data_o = 32'h00000000 /* 0x071c */;
                456: data_o = 32'h00000000 /* 0x0720 */;
                457: data_o = 32'h00000000 /* 0x0724 */;
                458: data_o = 32'h00000000 /* 0x0728 */;
                459: data_o = 32'h00000000 /* 0x072c */;
                460: data_o = 32'h00000000 /* 0x0730 */;
                461: data_o = 32'h00000000 /* 0x0734 */;
                462: data_o = 32'h00000000 /* 0x0738 */;
                463: data_o = 32'h00000000 /* 0x073c */;
                464: data_o = 32'h00000000 /* 0x0740 */;
                465: data_o = 32'h00000000 /* 0x0744 */;
                466: data_o = 32'h00000000 /* 0x0748 */;
                467: data_o = 32'h00000000 /* 0x074c */;
                468: data_o = 32'h00000000 /* 0x0750 */;
                469: data_o = 32'h00000000 /* 0x0754 */;
                470: data_o = 32'h00000000 /* 0x0758 */;
                471: data_o = 32'h00000000 /* 0x075c */;
                472: data_o = 32'h00000000 /* 0x0760 */;
                473: data_o = 32'h00000000 /* 0x0764 */;
                474: data_o = 32'h00000000 /* 0x0768 */;
                475: data_o = 32'h00000000 /* 0x076c */;
                476: data_o = 32'h00000000 /* 0x0770 */;
                477: data_o = 32'h00000000 /* 0x0774 */;
                478: data_o = 32'h00000000 /* 0x0778 */;
                479: data_o = 32'h00000000 /* 0x077c */;
                480: data_o = 32'h00000000 /* 0x0780 */;
                481: data_o = 32'h00000000 /* 0x0784 */;
                482: data_o = 32'h00000000 /* 0x0788 */;
                483: data_o = 32'h00000000 /* 0x078c */;
                484: data_o = 32'h00000000 /* 0x0790 */;
                485: data_o = 32'h00000000 /* 0x0794 */;
                486: data_o = 32'h00000000 /* 0x0798 */;
                487: data_o = 32'h00000000 /* 0x079c */;
                488: data_o = 32'h00000000 /* 0x07a0 */;
                489: data_o = 32'h00000000 /* 0x07a4 */;
                490: data_o = 32'h00000000 /* 0x07a8 */;
                491: data_o = 32'h00000000 /* 0x07ac */;
                492: data_o = 32'h00000000 /* 0x07b0 */;
                493: data_o = 32'h00000000 /* 0x07b4 */;
                494: data_o = 32'h00000000 /* 0x07b8 */;
                495: data_o = 32'h00000000 /* 0x07bc */;
                496: data_o = 32'h00000000 /* 0x07c0 */;
                497: data_o = 32'h00000000 /* 0x07c4 */;
                498: data_o = 32'h00000000 /* 0x07c8 */;
                499: data_o = 32'h00000000 /* 0x07cc */;
                500: data_o = 32'h00000000 /* 0x07d0 */;
                501: data_o = 32'h00000000 /* 0x07d4 */;
                502: data_o = 32'h00000000 /* 0x07d8 */;
                503: data_o = 32'h00000000 /* 0x07dc */;
                504: data_o = 32'h00000000 /* 0x07e0 */;
                505: data_o = 32'h00000000 /* 0x07e4 */;
                506: data_o = 32'h00000000 /* 0x07e8 */;
                507: data_o = 32'h00000000 /* 0x07ec */;
                508: data_o = 32'h00000000 /* 0x07f0 */;
                509: data_o = 32'h00000000 /* 0x07f4 */;
                510: data_o = 32'h00000000 /* 0x07f8 */;
                511: data_o = 32'h00000000 /* 0x07fc */;
                512: data_o = 32'h00000000 /* 0x0800 */;
                513: data_o = 32'h00000000 /* 0x0804 */;
                514: data_o = 32'h00000000 /* 0x0808 */;
                515: data_o = 32'h00000000 /* 0x080c */;
                516: data_o = 32'h00000000 /* 0x0810 */;
                517: data_o = 32'h00000000 /* 0x0814 */;
                518: data_o = 32'h00000000 /* 0x0818 */;
                519: data_o = 32'h00000000 /* 0x081c */;
                520: data_o = 32'h00000000 /* 0x0820 */;
                521: data_o = 32'h00000000 /* 0x0824 */;
                522: data_o = 32'h00000000 /* 0x0828 */;
                523: data_o = 32'h00000000 /* 0x082c */;
                524: data_o = 32'h00000000 /* 0x0830 */;
                525: data_o = 32'h00000000 /* 0x0834 */;
                526: data_o = 32'h00000000 /* 0x0838 */;
                527: data_o = 32'h00000000 /* 0x083c */;
                528: data_o = 32'h00000000 /* 0x0840 */;
                529: data_o = 32'h00000000 /* 0x0844 */;
                530: data_o = 32'h00000000 /* 0x0848 */;
                531: data_o = 32'h00000000 /* 0x084c */;
                532: data_o = 32'h00000000 /* 0x0850 */;
                533: data_o = 32'h00000000 /* 0x0854 */;
                534: data_o = 32'h00000000 /* 0x0858 */;
                535: data_o = 32'h00000000 /* 0x085c */;
                536: data_o = 32'h00000000 /* 0x0860 */;
                537: data_o = 32'h00000000 /* 0x0864 */;
                538: data_o = 32'h00000000 /* 0x0868 */;
                539: data_o = 32'h00000000 /* 0x086c */;
                540: data_o = 32'h00000000 /* 0x0870 */;
                541: data_o = 32'h00000000 /* 0x0874 */;
                542: data_o = 32'h00000000 /* 0x0878 */;
                543: data_o = 32'h00000000 /* 0x087c */;
                544: data_o = 32'h00000000 /* 0x0880 */;
                545: data_o = 32'h00000000 /* 0x0884 */;
                546: data_o = 32'h00000000 /* 0x0888 */;
                547: data_o = 32'h00000000 /* 0x088c */;
                548: data_o = 32'h00000000 /* 0x0890 */;
                549: data_o = 32'h00000000 /* 0x0894 */;
                550: data_o = 32'h00000000 /* 0x0898 */;
                551: data_o = 32'h00000000 /* 0x089c */;
                552: data_o = 32'h00000000 /* 0x08a0 */;
                553: data_o = 32'h00000000 /* 0x08a4 */;
                554: data_o = 32'h00000000 /* 0x08a8 */;
                555: data_o = 32'h00000000 /* 0x08ac */;
                556: data_o = 32'h00000000 /* 0x08b0 */;
                557: data_o = 32'h00000000 /* 0x08b4 */;
                558: data_o = 32'h00000000 /* 0x08b8 */;
                559: data_o = 32'h00000000 /* 0x08bc */;
                560: data_o = 32'h00000000 /* 0x08c0 */;
                561: data_o = 32'h00000000 /* 0x08c4 */;
                562: data_o = 32'h00000000 /* 0x08c8 */;
                563: data_o = 32'h00000000 /* 0x08cc */;
                564: data_o = 32'h00000000 /* 0x08d0 */;
                565: data_o = 32'h00000000 /* 0x08d4 */;
                566: data_o = 32'h00000000 /* 0x08d8 */;
                567: data_o = 32'h00000000 /* 0x08dc */;
                568: data_o = 32'h00000000 /* 0x08e0 */;
                569: data_o = 32'h00000000 /* 0x08e4 */;
                570: data_o = 32'h00000000 /* 0x08e8 */;
                571: data_o = 32'h00000000 /* 0x08ec */;
                572: data_o = 32'h00000000 /* 0x08f0 */;
                573: data_o = 32'h00000000 /* 0x08f4 */;
                574: data_o = 32'h00000000 /* 0x08f8 */;
                575: data_o = 32'h00000000 /* 0x08fc */;
                576: data_o = 32'h00000000 /* 0x0900 */;
                577: data_o = 32'h00000000 /* 0x0904 */;
                578: data_o = 32'h00000000 /* 0x0908 */;
                579: data_o = 32'h00000000 /* 0x090c */;
                580: data_o = 32'h00000000 /* 0x0910 */;
                581: data_o = 32'h00000000 /* 0x0914 */;
                582: data_o = 32'h00000000 /* 0x0918 */;
                583: data_o = 32'h00000000 /* 0x091c */;
                584: data_o = 32'h00000000 /* 0x0920 */;
                585: data_o = 32'h00000000 /* 0x0924 */;
                586: data_o = 32'h00000000 /* 0x0928 */;
                587: data_o = 32'h00000000 /* 0x092c */;
                588: data_o = 32'h00000000 /* 0x0930 */;
                589: data_o = 32'h00000000 /* 0x0934 */;
                590: data_o = 32'h00000000 /* 0x0938 */;
                591: data_o = 32'h00000000 /* 0x093c */;
                592: data_o = 32'h00000000 /* 0x0940 */;
                593: data_o = 32'h00000000 /* 0x0944 */;
                594: data_o = 32'h00000000 /* 0x0948 */;
                595: data_o = 32'h00000000 /* 0x094c */;
                596: data_o = 32'h00000000 /* 0x0950 */;
                597: data_o = 32'h00000000 /* 0x0954 */;
                598: data_o = 32'h00000000 /* 0x0958 */;
                599: data_o = 32'h00000000 /* 0x095c */;
                600: data_o = 32'h00000000 /* 0x0960 */;
                601: data_o = 32'h00000000 /* 0x0964 */;
                602: data_o = 32'h00000000 /* 0x0968 */;
                603: data_o = 32'h00000000 /* 0x096c */;
                604: data_o = 32'h00000000 /* 0x0970 */;
                605: data_o = 32'h00000000 /* 0x0974 */;
                606: data_o = 32'h00000000 /* 0x0978 */;
                607: data_o = 32'h00000000 /* 0x097c */;
                608: data_o = 32'h00000000 /* 0x0980 */;
                609: data_o = 32'h00000000 /* 0x0984 */;
                610: data_o = 32'h00000000 /* 0x0988 */;
                611: data_o = 32'h00000000 /* 0x098c */;
                612: data_o = 32'h00000000 /* 0x0990 */;
                613: data_o = 32'h00000000 /* 0x0994 */;
                614: data_o = 32'h00000000 /* 0x0998 */;
                615: data_o = 32'h00000000 /* 0x099c */;
                616: data_o = 32'h00000000 /* 0x09a0 */;
                617: data_o = 32'h00000000 /* 0x09a4 */;
                618: data_o = 32'h00000000 /* 0x09a8 */;
                619: data_o = 32'h00000000 /* 0x09ac */;
                620: data_o = 32'h00000000 /* 0x09b0 */;
                621: data_o = 32'h00000000 /* 0x09b4 */;
                622: data_o = 32'h00000000 /* 0x09b8 */;
                623: data_o = 32'h00000000 /* 0x09bc */;
                624: data_o = 32'h00000000 /* 0x09c0 */;
                625: data_o = 32'h00000000 /* 0x09c4 */;
                626: data_o = 32'h00000000 /* 0x09c8 */;
                627: data_o = 32'h00000000 /* 0x09cc */;
                628: data_o = 32'h00000000 /* 0x09d0 */;
                629: data_o = 32'h00000000 /* 0x09d4 */;
                630: data_o = 32'h00000000 /* 0x09d8 */;
                631: data_o = 32'h00000000 /* 0x09dc */;
                632: data_o = 32'h00000000 /* 0x09e0 */;
                633: data_o = 32'h00000000 /* 0x09e4 */;
                634: data_o = 32'h00000000 /* 0x09e8 */;
                635: data_o = 32'h00000000 /* 0x09ec */;
                636: data_o = 32'h00000000 /* 0x09f0 */;
                637: data_o = 32'h00000000 /* 0x09f4 */;
                638: data_o = 32'h00000000 /* 0x09f8 */;
                639: data_o = 32'h00000000 /* 0x09fc */;
                640: data_o = 32'h00000000 /* 0x0a00 */;
                641: data_o = 32'h00000000 /* 0x0a04 */;
                642: data_o = 32'h00000000 /* 0x0a08 */;
                643: data_o = 32'h00000000 /* 0x0a0c */;
                644: data_o = 32'h00000000 /* 0x0a10 */;
                645: data_o = 32'h00000000 /* 0x0a14 */;
                646: data_o = 32'h00000000 /* 0x0a18 */;
                647: data_o = 32'h00000000 /* 0x0a1c */;
                648: data_o = 32'h00000000 /* 0x0a20 */;
                649: data_o = 32'h00000000 /* 0x0a24 */;
                650: data_o = 32'h00000000 /* 0x0a28 */;
                651: data_o = 32'h00000000 /* 0x0a2c */;
                652: data_o = 32'h00000000 /* 0x0a30 */;
                653: data_o = 32'h00000000 /* 0x0a34 */;
                654: data_o = 32'h00000000 /* 0x0a38 */;
                655: data_o = 32'h00000000 /* 0x0a3c */;
                656: data_o = 32'h00000000 /* 0x0a40 */;
                657: data_o = 32'h00000000 /* 0x0a44 */;
                658: data_o = 32'h00000000 /* 0x0a48 */;
                659: data_o = 32'h00000000 /* 0x0a4c */;
                660: data_o = 32'h00000000 /* 0x0a50 */;
                661: data_o = 32'h00000000 /* 0x0a54 */;
                662: data_o = 32'h00000000 /* 0x0a58 */;
                663: data_o = 32'h00000000 /* 0x0a5c */;
                664: data_o = 32'h00000000 /* 0x0a60 */;
                665: data_o = 32'h00000000 /* 0x0a64 */;
                666: data_o = 32'h00000000 /* 0x0a68 */;
                667: data_o = 32'h00000000 /* 0x0a6c */;
                668: data_o = 32'h00000000 /* 0x0a70 */;
                669: data_o = 32'h00000000 /* 0x0a74 */;
                670: data_o = 32'h00000000 /* 0x0a78 */;
                671: data_o = 32'h00000000 /* 0x0a7c */;
                672: data_o = 32'h00000000 /* 0x0a80 */;
                673: data_o = 32'h00000000 /* 0x0a84 */;
                674: data_o = 32'h00000000 /* 0x0a88 */;
                675: data_o = 32'h00000000 /* 0x0a8c */;
                676: data_o = 32'h00000000 /* 0x0a90 */;
                677: data_o = 32'h00000000 /* 0x0a94 */;
                678: data_o = 32'h00000000 /* 0x0a98 */;
                679: data_o = 32'h00000000 /* 0x0a9c */;
                680: data_o = 32'h00000000 /* 0x0aa0 */;
                681: data_o = 32'h00000000 /* 0x0aa4 */;
                682: data_o = 32'h00000000 /* 0x0aa8 */;
                683: data_o = 32'h00000000 /* 0x0aac */;
                684: data_o = 32'h00000000 /* 0x0ab0 */;
                685: data_o = 32'h00000000 /* 0x0ab4 */;
                686: data_o = 32'h00000000 /* 0x0ab8 */;
                687: data_o = 32'h00000000 /* 0x0abc */;
                688: data_o = 32'h00000000 /* 0x0ac0 */;
                689: data_o = 32'h00000000 /* 0x0ac4 */;
                690: data_o = 32'h00000000 /* 0x0ac8 */;
                691: data_o = 32'h00000000 /* 0x0acc */;
                692: data_o = 32'h00000000 /* 0x0ad0 */;
                693: data_o = 32'h00000000 /* 0x0ad4 */;
                694: data_o = 32'h00000000 /* 0x0ad8 */;
                695: data_o = 32'h00000000 /* 0x0adc */;
                696: data_o = 32'h00000000 /* 0x0ae0 */;
                697: data_o = 32'h00000000 /* 0x0ae4 */;
                698: data_o = 32'h00000000 /* 0x0ae8 */;
                699: data_o = 32'h00000000 /* 0x0aec */;
                700: data_o = 32'h00000000 /* 0x0af0 */;
                701: data_o = 32'h00000000 /* 0x0af4 */;
                702: data_o = 32'h00000000 /* 0x0af8 */;
                703: data_o = 32'h00000000 /* 0x0afc */;
                704: data_o = 32'h00000000 /* 0x0b00 */;
                705: data_o = 32'h00000000 /* 0x0b04 */;
                706: data_o = 32'h00000000 /* 0x0b08 */;
                707: data_o = 32'h00000000 /* 0x0b0c */;
                708: data_o = 32'h00000000 /* 0x0b10 */;
                709: data_o = 32'h00000000 /* 0x0b14 */;
                710: data_o = 32'h00000000 /* 0x0b18 */;
                711: data_o = 32'h00000000 /* 0x0b1c */;
                712: data_o = 32'h00000000 /* 0x0b20 */;
                713: data_o = 32'h00000000 /* 0x0b24 */;
                714: data_o = 32'h00000000 /* 0x0b28 */;
                715: data_o = 32'h00000000 /* 0x0b2c */;
                716: data_o = 32'h00000000 /* 0x0b30 */;
                717: data_o = 32'h00000000 /* 0x0b34 */;
                718: data_o = 32'h00000000 /* 0x0b38 */;
                719: data_o = 32'h00000000 /* 0x0b3c */;
                720: data_o = 32'h00000000 /* 0x0b40 */;
                721: data_o = 32'h00000000 /* 0x0b44 */;
                722: data_o = 32'h00000000 /* 0x0b48 */;
                723: data_o = 32'h00000000 /* 0x0b4c */;
                724: data_o = 32'h00000000 /* 0x0b50 */;
                725: data_o = 32'h00000000 /* 0x0b54 */;
                726: data_o = 32'h00000000 /* 0x0b58 */;
                727: data_o = 32'h00000000 /* 0x0b5c */;
                728: data_o = 32'h00000000 /* 0x0b60 */;
                729: data_o = 32'h00000000 /* 0x0b64 */;
                730: data_o = 32'h00000000 /* 0x0b68 */;
                731: data_o = 32'h00000000 /* 0x0b6c */;
                732: data_o = 32'h00000000 /* 0x0b70 */;
                733: data_o = 32'h00000000 /* 0x0b74 */;
                734: data_o = 32'h00000000 /* 0x0b78 */;
                735: data_o = 32'h00000000 /* 0x0b7c */;
                736: data_o = 32'h00000000 /* 0x0b80 */;
                737: data_o = 32'h00000000 /* 0x0b84 */;
                738: data_o = 32'h00000000 /* 0x0b88 */;
                739: data_o = 32'h00000000 /* 0x0b8c */;
                740: data_o = 32'h00000000 /* 0x0b90 */;
                741: data_o = 32'h00000000 /* 0x0b94 */;
                742: data_o = 32'h00000000 /* 0x0b98 */;
                743: data_o = 32'h00000000 /* 0x0b9c */;
                744: data_o = 32'h00000000 /* 0x0ba0 */;
                745: data_o = 32'h00000000 /* 0x0ba4 */;
                746: data_o = 32'h00000000 /* 0x0ba8 */;
                747: data_o = 32'h00000000 /* 0x0bac */;
                748: data_o = 32'h00000000 /* 0x0bb0 */;
                749: data_o = 32'h00000000 /* 0x0bb4 */;
                750: data_o = 32'h00000000 /* 0x0bb8 */;
                751: data_o = 32'h00000000 /* 0x0bbc */;
                752: data_o = 32'h00000000 /* 0x0bc0 */;
                753: data_o = 32'h00000000 /* 0x0bc4 */;
                754: data_o = 32'h00000000 /* 0x0bc8 */;
                755: data_o = 32'h00000000 /* 0x0bcc */;
                756: data_o = 32'h00000000 /* 0x0bd0 */;
                757: data_o = 32'h00000000 /* 0x0bd4 */;
                758: data_o = 32'h00000000 /* 0x0bd8 */;
                759: data_o = 32'h00000000 /* 0x0bdc */;
                760: data_o = 32'h00000000 /* 0x0be0 */;
                761: data_o = 32'h00000000 /* 0x0be4 */;
                762: data_o = 32'h00000000 /* 0x0be8 */;
                763: data_o = 32'h00000000 /* 0x0bec */;
                764: data_o = 32'h00000000 /* 0x0bf0 */;
                765: data_o = 32'h00000000 /* 0x0bf4 */;
                766: data_o = 32'h00000000 /* 0x0bf8 */;
                767: data_o = 32'h00000000 /* 0x0bfc */;
                768: data_o = 32'h00000000 /* 0x0c00 */;
                769: data_o = 32'h00000000 /* 0x0c04 */;
                770: data_o = 32'h00000000 /* 0x0c08 */;
                771: data_o = 32'h00000000 /* 0x0c0c */;
                772: data_o = 32'h00000000 /* 0x0c10 */;
                773: data_o = 32'h00000000 /* 0x0c14 */;
                774: data_o = 32'h00000000 /* 0x0c18 */;
                775: data_o = 32'h00000000 /* 0x0c1c */;
                776: data_o = 32'h00000000 /* 0x0c20 */;
                777: data_o = 32'h00000000 /* 0x0c24 */;
                778: data_o = 32'h00000000 /* 0x0c28 */;
                779: data_o = 32'h00000000 /* 0x0c2c */;
                780: data_o = 32'h00000000 /* 0x0c30 */;
                781: data_o = 32'h00000000 /* 0x0c34 */;
                782: data_o = 32'h00000000 /* 0x0c38 */;
                783: data_o = 32'h00000000 /* 0x0c3c */;
                784: data_o = 32'h00000000 /* 0x0c40 */;
                785: data_o = 32'h00000000 /* 0x0c44 */;
                786: data_o = 32'h00000000 /* 0x0c48 */;
                787: data_o = 32'h00000000 /* 0x0c4c */;
                788: data_o = 32'h00000000 /* 0x0c50 */;
                789: data_o = 32'h00000000 /* 0x0c54 */;
                790: data_o = 32'h00000000 /* 0x0c58 */;
                791: data_o = 32'h00000000 /* 0x0c5c */;
                792: data_o = 32'h00000000 /* 0x0c60 */;
                793: data_o = 32'h00000000 /* 0x0c64 */;
                794: data_o = 32'h00000000 /* 0x0c68 */;
                795: data_o = 32'h00000000 /* 0x0c6c */;
                796: data_o = 32'h00000000 /* 0x0c70 */;
                797: data_o = 32'h00000000 /* 0x0c74 */;
                798: data_o = 32'h00000000 /* 0x0c78 */;
                799: data_o = 32'h00000000 /* 0x0c7c */;
                800: data_o = 32'h00000000 /* 0x0c80 */;
                801: data_o = 32'h00000000 /* 0x0c84 */;
                802: data_o = 32'h00000000 /* 0x0c88 */;
                803: data_o = 32'h00000000 /* 0x0c8c */;
                804: data_o = 32'h00000000 /* 0x0c90 */;
                805: data_o = 32'h00000000 /* 0x0c94 */;
                806: data_o = 32'h00000000 /* 0x0c98 */;
                807: data_o = 32'h00000000 /* 0x0c9c */;
                808: data_o = 32'h00000000 /* 0x0ca0 */;
                809: data_o = 32'h00000000 /* 0x0ca4 */;
                810: data_o = 32'h00000000 /* 0x0ca8 */;
                811: data_o = 32'h00000000 /* 0x0cac */;
                812: data_o = 32'h00000000 /* 0x0cb0 */;
                813: data_o = 32'h00000000 /* 0x0cb4 */;
                814: data_o = 32'h00000000 /* 0x0cb8 */;
                815: data_o = 32'h00000000 /* 0x0cbc */;
                816: data_o = 32'h00000000 /* 0x0cc0 */;
                817: data_o = 32'h00000000 /* 0x0cc4 */;
                818: data_o = 32'h00000000 /* 0x0cc8 */;
                819: data_o = 32'h00000000 /* 0x0ccc */;
                820: data_o = 32'h00000000 /* 0x0cd0 */;
                821: data_o = 32'h00000000 /* 0x0cd4 */;
                822: data_o = 32'h00000000 /* 0x0cd8 */;
                823: data_o = 32'h00000000 /* 0x0cdc */;
                824: data_o = 32'h00000000 /* 0x0ce0 */;
                825: data_o = 32'h00000000 /* 0x0ce4 */;
                826: data_o = 32'h00000000 /* 0x0ce8 */;
                827: data_o = 32'h00000000 /* 0x0cec */;
                828: data_o = 32'h00000000 /* 0x0cf0 */;
                829: data_o = 32'h00000000 /* 0x0cf4 */;
                830: data_o = 32'h00000000 /* 0x0cf8 */;
                831: data_o = 32'h00000000 /* 0x0cfc */;
                832: data_o = 32'h00000000 /* 0x0d00 */;
                833: data_o = 32'h00000000 /* 0x0d04 */;
                834: data_o = 32'h00000000 /* 0x0d08 */;
                835: data_o = 32'h00000000 /* 0x0d0c */;
                836: data_o = 32'h00000000 /* 0x0d10 */;
                837: data_o = 32'h00000000 /* 0x0d14 */;
                838: data_o = 32'h00000000 /* 0x0d18 */;
                839: data_o = 32'h00000000 /* 0x0d1c */;
                840: data_o = 32'h00000000 /* 0x0d20 */;
                841: data_o = 32'h00000000 /* 0x0d24 */;
                842: data_o = 32'h00000000 /* 0x0d28 */;
                843: data_o = 32'h00000000 /* 0x0d2c */;
                844: data_o = 32'h00000000 /* 0x0d30 */;
                845: data_o = 32'h00000000 /* 0x0d34 */;
                846: data_o = 32'h00000000 /* 0x0d38 */;
                847: data_o = 32'h00000000 /* 0x0d3c */;
                848: data_o = 32'h00000000 /* 0x0d40 */;
                849: data_o = 32'h00000000 /* 0x0d44 */;
                850: data_o = 32'h00000000 /* 0x0d48 */;
                851: data_o = 32'h00000000 /* 0x0d4c */;
                852: data_o = 32'h00000000 /* 0x0d50 */;
                853: data_o = 32'h00000000 /* 0x0d54 */;
                854: data_o = 32'h00000000 /* 0x0d58 */;
                855: data_o = 32'h00000000 /* 0x0d5c */;
                856: data_o = 32'h00000000 /* 0x0d60 */;
                857: data_o = 32'h00000000 /* 0x0d64 */;
                858: data_o = 32'h00000000 /* 0x0d68 */;
                859: data_o = 32'h00000000 /* 0x0d6c */;
                860: data_o = 32'h00000000 /* 0x0d70 */;
                861: data_o = 32'h00000000 /* 0x0d74 */;
                862: data_o = 32'h00000000 /* 0x0d78 */;
                863: data_o = 32'h00000000 /* 0x0d7c */;
                864: data_o = 32'h00000000 /* 0x0d80 */;
                865: data_o = 32'h00000000 /* 0x0d84 */;
                866: data_o = 32'h00000000 /* 0x0d88 */;
                867: data_o = 32'h00000000 /* 0x0d8c */;
                868: data_o = 32'h00000000 /* 0x0d90 */;
                869: data_o = 32'h00000000 /* 0x0d94 */;
                870: data_o = 32'h00000000 /* 0x0d98 */;
                871: data_o = 32'h00000000 /* 0x0d9c */;
                872: data_o = 32'h00000000 /* 0x0da0 */;
                873: data_o = 32'h00000000 /* 0x0da4 */;
                874: data_o = 32'h00000000 /* 0x0da8 */;
                875: data_o = 32'h00000000 /* 0x0dac */;
                876: data_o = 32'h00000000 /* 0x0db0 */;
                877: data_o = 32'h00000000 /* 0x0db4 */;
                878: data_o = 32'h00000000 /* 0x0db8 */;
                879: data_o = 32'h00000000 /* 0x0dbc */;
                880: data_o = 32'h00000000 /* 0x0dc0 */;
                881: data_o = 32'h00000000 /* 0x0dc4 */;
                882: data_o = 32'h00000000 /* 0x0dc8 */;
                883: data_o = 32'h00000000 /* 0x0dcc */;
                884: data_o = 32'h00000000 /* 0x0dd0 */;
                885: data_o = 32'h00000000 /* 0x0dd4 */;
                886: data_o = 32'h00000000 /* 0x0dd8 */;
                887: data_o = 32'h00000000 /* 0x0ddc */;
                888: data_o = 32'h00000000 /* 0x0de0 */;
                889: data_o = 32'h00000000 /* 0x0de4 */;
                890: data_o = 32'h00000000 /* 0x0de8 */;
                891: data_o = 32'h00000000 /* 0x0dec */;
                892: data_o = 32'h00000000 /* 0x0df0 */;
                893: data_o = 32'h00000000 /* 0x0df4 */;
                894: data_o = 32'h00000000 /* 0x0df8 */;
                895: data_o = 32'h00000000 /* 0x0dfc */;
                896: data_o = 32'h00000000 /* 0x0e00 */;
                897: data_o = 32'h00000000 /* 0x0e04 */;
                898: data_o = 32'h00000000 /* 0x0e08 */;
                899: data_o = 32'h00000000 /* 0x0e0c */;
                900: data_o = 32'h00000000 /* 0x0e10 */;
                901: data_o = 32'h00000000 /* 0x0e14 */;
                902: data_o = 32'h00000000 /* 0x0e18 */;
                903: data_o = 32'h00000000 /* 0x0e1c */;
                904: data_o = 32'h00000000 /* 0x0e20 */;
                905: data_o = 32'h00000000 /* 0x0e24 */;
                906: data_o = 32'h00000000 /* 0x0e28 */;
                907: data_o = 32'h00000000 /* 0x0e2c */;
                908: data_o = 32'h00000000 /* 0x0e30 */;
                909: data_o = 32'h00000000 /* 0x0e34 */;
                910: data_o = 32'h00000000 /* 0x0e38 */;
                911: data_o = 32'h00000000 /* 0x0e3c */;
                912: data_o = 32'h00000000 /* 0x0e40 */;
                913: data_o = 32'h00000000 /* 0x0e44 */;
                914: data_o = 32'h00000000 /* 0x0e48 */;
                915: data_o = 32'h00000000 /* 0x0e4c */;
                916: data_o = 32'h00000000 /* 0x0e50 */;
                917: data_o = 32'h00000000 /* 0x0e54 */;
                918: data_o = 32'h00000000 /* 0x0e58 */;
                919: data_o = 32'h00000000 /* 0x0e5c */;
                920: data_o = 32'h00000000 /* 0x0e60 */;
                921: data_o = 32'h00000000 /* 0x0e64 */;
                922: data_o = 32'h00000000 /* 0x0e68 */;
                923: data_o = 32'h00000000 /* 0x0e6c */;
                924: data_o = 32'h00000000 /* 0x0e70 */;
                925: data_o = 32'h00000000 /* 0x0e74 */;
                926: data_o = 32'h00000000 /* 0x0e78 */;
                927: data_o = 32'h00000000 /* 0x0e7c */;
                928: data_o = 32'h00000000 /* 0x0e80 */;
                929: data_o = 32'h00000000 /* 0x0e84 */;
                930: data_o = 32'h00000000 /* 0x0e88 */;
                931: data_o = 32'h00000000 /* 0x0e8c */;
                932: data_o = 32'h00000000 /* 0x0e90 */;
                933: data_o = 32'h00000000 /* 0x0e94 */;
                934: data_o = 32'h00000000 /* 0x0e98 */;
                935: data_o = 32'h00000000 /* 0x0e9c */;
                936: data_o = 32'h00000000 /* 0x0ea0 */;
                937: data_o = 32'h00000000 /* 0x0ea4 */;
                938: data_o = 32'h00000000 /* 0x0ea8 */;
                939: data_o = 32'h00000000 /* 0x0eac */;
                940: data_o = 32'h00000000 /* 0x0eb0 */;
                941: data_o = 32'h00000000 /* 0x0eb4 */;
                942: data_o = 32'h00000000 /* 0x0eb8 */;
                943: data_o = 32'h00000000 /* 0x0ebc */;
                944: data_o = 32'h00000000 /* 0x0ec0 */;
                945: data_o = 32'h00000000 /* 0x0ec4 */;
                946: data_o = 32'h00000000 /* 0x0ec8 */;
                947: data_o = 32'h00000000 /* 0x0ecc */;
                948: data_o = 32'h00000000 /* 0x0ed0 */;
                949: data_o = 32'h00000000 /* 0x0ed4 */;
                950: data_o = 32'h00000000 /* 0x0ed8 */;
                951: data_o = 32'h00000000 /* 0x0edc */;
                952: data_o = 32'h00000000 /* 0x0ee0 */;
                953: data_o = 32'h00000000 /* 0x0ee4 */;
                954: data_o = 32'h00000000 /* 0x0ee8 */;
                955: data_o = 32'h00000000 /* 0x0eec */;
                956: data_o = 32'h00000000 /* 0x0ef0 */;
                957: data_o = 32'h00000000 /* 0x0ef4 */;
                958: data_o = 32'h00000000 /* 0x0ef8 */;
                959: data_o = 32'h00000000 /* 0x0efc */;
                960: data_o = 32'h00000000 /* 0x0f00 */;
                961: data_o = 32'h00000000 /* 0x0f04 */;
                962: data_o = 32'h00000000 /* 0x0f08 */;
                963: data_o = 32'h00000000 /* 0x0f0c */;
                964: data_o = 32'h00000000 /* 0x0f10 */;
                965: data_o = 32'h00000000 /* 0x0f14 */;
                966: data_o = 32'h00000000 /* 0x0f18 */;
                967: data_o = 32'h00000000 /* 0x0f1c */;
                968: data_o = 32'h00000000 /* 0x0f20 */;
                969: data_o = 32'h00000000 /* 0x0f24 */;
                970: data_o = 32'h00000000 /* 0x0f28 */;
                971: data_o = 32'h00000000 /* 0x0f2c */;
                972: data_o = 32'h00000000 /* 0x0f30 */;
                973: data_o = 32'h00000000 /* 0x0f34 */;
                974: data_o = 32'h00000000 /* 0x0f38 */;
                975: data_o = 32'h00000000 /* 0x0f3c */;
                976: data_o = 32'h00000000 /* 0x0f40 */;
                977: data_o = 32'h00000000 /* 0x0f44 */;
                978: data_o = 32'h00000000 /* 0x0f48 */;
                979: data_o = 32'h00000000 /* 0x0f4c */;
                980: data_o = 32'h00000000 /* 0x0f50 */;
                981: data_o = 32'h00000000 /* 0x0f54 */;
                982: data_o = 32'h00000000 /* 0x0f58 */;
                983: data_o = 32'h00000000 /* 0x0f5c */;
                984: data_o = 32'h00000000 /* 0x0f60 */;
                985: data_o = 32'h00000000 /* 0x0f64 */;
                986: data_o = 32'h00000000 /* 0x0f68 */;
                987: data_o = 32'h00000000 /* 0x0f6c */;
                988: data_o = 32'h00000000 /* 0x0f70 */;
                989: data_o = 32'h00000000 /* 0x0f74 */;
                990: data_o = 32'h00000000 /* 0x0f78 */;
                991: data_o = 32'h00000000 /* 0x0f7c */;
                992: data_o = 32'h00000000 /* 0x0f80 */;
                993: data_o = 32'h00000000 /* 0x0f84 */;
                994: data_o = 32'h00000000 /* 0x0f88 */;
                995: data_o = 32'h00000000 /* 0x0f8c */;
                996: data_o = 32'h00000000 /* 0x0f90 */;
                997: data_o = 32'h00000000 /* 0x0f94 */;
                998: data_o = 32'h00000000 /* 0x0f98 */;
                999: data_o = 32'h00000000 /* 0x0f9c */;
                1000: data_o = 32'h00000000 /* 0x0fa0 */;
                1001: data_o = 32'h00000000 /* 0x0fa4 */;
                1002: data_o = 32'h00000000 /* 0x0fa8 */;
                1003: data_o = 32'h00000000 /* 0x0fac */;
                1004: data_o = 32'h00000000 /* 0x0fb0 */;
                1005: data_o = 32'h00000000 /* 0x0fb4 */;
                1006: data_o = 32'h00000000 /* 0x0fb8 */;
                1007: data_o = 32'h00000000 /* 0x0fbc */;
                1008: data_o = 32'h00000000 /* 0x0fc0 */;
                1009: data_o = 32'h00000000 /* 0x0fc4 */;
                1010: data_o = 32'h00000000 /* 0x0fc8 */;
                1011: data_o = 32'h00000000 /* 0x0fcc */;
                1012: data_o = 32'h00000000 /* 0x0fd0 */;
                1013: data_o = 32'h00000000 /* 0x0fd4 */;
                1014: data_o = 32'h00000000 /* 0x0fd8 */;
                1015: data_o = 32'h00000000 /* 0x0fdc */;
                1016: data_o = 32'h00000000 /* 0x0fe0 */;
                1017: data_o = 32'h00000000 /* 0x0fe4 */;
                1018: data_o = 32'h00000000 /* 0x0fe8 */;
                1019: data_o = 32'h00000000 /* 0x0fec */;
                1020: data_o = 32'h00000000 /* 0x0ff0 */;
                1021: data_o = 32'h00000000 /* 0x0ff4 */;
                1022: data_o = 32'h00000000 /* 0x0ff8 */;
                1023: data_o = 32'h00000000 /* 0x0ffc */;
                1024: data_o = 32'h00000000 /* 0x1000 */;
                1025: data_o = 32'h00000000 /* 0x1004 */;
                1026: data_o = 32'h00000000 /* 0x1008 */;
                1027: data_o = 32'h00000000 /* 0x100c */;
                1028: data_o = 32'h00000000 /* 0x1010 */;
                1029: data_o = 32'h00000000 /* 0x1014 */;
                1030: data_o = 32'h00000000 /* 0x1018 */;
                1031: data_o = 32'h00000000 /* 0x101c */;
                1032: data_o = 32'h00000000 /* 0x1020 */;
                1033: data_o = 32'h00000000 /* 0x1024 */;
                1034: data_o = 32'h00000000 /* 0x1028 */;
                1035: data_o = 32'h00000000 /* 0x102c */;
                1036: data_o = 32'h00000000 /* 0x1030 */;
                1037: data_o = 32'h00000000 /* 0x1034 */;
                1038: data_o = 32'h00000000 /* 0x1038 */;
                1039: data_o = 32'h00000000 /* 0x103c */;
                1040: data_o = 32'h00000000 /* 0x1040 */;
                1041: data_o = 32'h00000000 /* 0x1044 */;
                1042: data_o = 32'h00000000 /* 0x1048 */;
                1043: data_o = 32'h00000000 /* 0x104c */;
                1044: data_o = 32'h00000000 /* 0x1050 */;
                1045: data_o = 32'h00000000 /* 0x1054 */;
                1046: data_o = 32'h00000000 /* 0x1058 */;
                1047: data_o = 32'h00000000 /* 0x105c */;
                1048: data_o = 32'h00000000 /* 0x1060 */;
                1049: data_o = 32'h00000000 /* 0x1064 */;
                1050: data_o = 32'h00000000 /* 0x1068 */;
                1051: data_o = 32'h00000000 /* 0x106c */;
                1052: data_o = 32'h00000000 /* 0x1070 */;
                1053: data_o = 32'h00000000 /* 0x1074 */;
                1054: data_o = 32'h00000000 /* 0x1078 */;
                1055: data_o = 32'h00000000 /* 0x107c */;
                1056: data_o = 32'h00000000 /* 0x1080 */;
                1057: data_o = 32'h00000000 /* 0x1084 */;
                1058: data_o = 32'h00000000 /* 0x1088 */;
                1059: data_o = 32'h00000000 /* 0x108c */;
                1060: data_o = 32'h00000000 /* 0x1090 */;
                1061: data_o = 32'h00000000 /* 0x1094 */;
                1062: data_o = 32'h00000000 /* 0x1098 */;
                1063: data_o = 32'h00000000 /* 0x109c */;
                1064: data_o = 32'h00000000 /* 0x10a0 */;
                1065: data_o = 32'h00000000 /* 0x10a4 */;
                1066: data_o = 32'h00000000 /* 0x10a8 */;
                1067: data_o = 32'h00000000 /* 0x10ac */;
                1068: data_o = 32'h00000000 /* 0x10b0 */;
                1069: data_o = 32'h00000000 /* 0x10b4 */;
                1070: data_o = 32'h00000000 /* 0x10b8 */;
                1071: data_o = 32'h00000000 /* 0x10bc */;
                1072: data_o = 32'h00000000 /* 0x10c0 */;
                1073: data_o = 32'h00000000 /* 0x10c4 */;
                1074: data_o = 32'h00000000 /* 0x10c8 */;
                1075: data_o = 32'h00000000 /* 0x10cc */;
                1076: data_o = 32'h00000000 /* 0x10d0 */;
                1077: data_o = 32'h00000000 /* 0x10d4 */;
                1078: data_o = 32'h00000000 /* 0x10d8 */;
                1079: data_o = 32'h00000000 /* 0x10dc */;
                1080: data_o = 32'h00000000 /* 0x10e0 */;
                1081: data_o = 32'h00000000 /* 0x10e4 */;
                1082: data_o = 32'h00000000 /* 0x10e8 */;
                1083: data_o = 32'h00000000 /* 0x10ec */;
                1084: data_o = 32'h00000000 /* 0x10f0 */;
                1085: data_o = 32'h00000000 /* 0x10f4 */;
                1086: data_o = 32'h00000000 /* 0x10f8 */;
                1087: data_o = 32'h00000000 /* 0x10fc */;
                1088: data_o = 32'h00000000 /* 0x1100 */;
                1089: data_o = 32'h00000000 /* 0x1104 */;
                1090: data_o = 32'h00000000 /* 0x1108 */;
                1091: data_o = 32'h00000000 /* 0x110c */;
                1092: data_o = 32'h00000000 /* 0x1110 */;
                1093: data_o = 32'h00000000 /* 0x1114 */;
                1094: data_o = 32'h00000000 /* 0x1118 */;
                1095: data_o = 32'h00000000 /* 0x111c */;
                1096: data_o = 32'h00000000 /* 0x1120 */;
                1097: data_o = 32'h00000000 /* 0x1124 */;
                1098: data_o = 32'h00000000 /* 0x1128 */;
                1099: data_o = 32'h00000000 /* 0x112c */;
                1100: data_o = 32'h00000000 /* 0x1130 */;
                1101: data_o = 32'h00000000 /* 0x1134 */;
                1102: data_o = 32'h00000000 /* 0x1138 */;
                1103: data_o = 32'h00000000 /* 0x113c */;
                1104: data_o = 32'h00000000 /* 0x1140 */;
                1105: data_o = 32'h00000000 /* 0x1144 */;
                1106: data_o = 32'h00000000 /* 0x1148 */;
                1107: data_o = 32'h00000000 /* 0x114c */;
                1108: data_o = 32'h00000000 /* 0x1150 */;
                1109: data_o = 32'h00000000 /* 0x1154 */;
                1110: data_o = 32'h00000000 /* 0x1158 */;
                1111: data_o = 32'h00000000 /* 0x115c */;
                1112: data_o = 32'h00000000 /* 0x1160 */;
                1113: data_o = 32'h00000000 /* 0x1164 */;
                1114: data_o = 32'h00000000 /* 0x1168 */;
                1115: data_o = 32'h00000000 /* 0x116c */;
                1116: data_o = 32'h00000000 /* 0x1170 */;
                1117: data_o = 32'h00000000 /* 0x1174 */;
                1118: data_o = 32'h00000000 /* 0x1178 */;
                1119: data_o = 32'h00000000 /* 0x117c */;
                1120: data_o = 32'h00000000 /* 0x1180 */;
                1121: data_o = 32'h00000000 /* 0x1184 */;
                1122: data_o = 32'h00000000 /* 0x1188 */;
                1123: data_o = 32'h00000000 /* 0x118c */;
                1124: data_o = 32'h00000000 /* 0x1190 */;
                1125: data_o = 32'h00000000 /* 0x1194 */;
                1126: data_o = 32'h00000000 /* 0x1198 */;
                1127: data_o = 32'h00000000 /* 0x119c */;
                1128: data_o = 32'h00000000 /* 0x11a0 */;
                1129: data_o = 32'h00000000 /* 0x11a4 */;
                1130: data_o = 32'h00000000 /* 0x11a8 */;
                1131: data_o = 32'h00000000 /* 0x11ac */;
                1132: data_o = 32'h00000000 /* 0x11b0 */;
                1133: data_o = 32'h00000000 /* 0x11b4 */;
                1134: data_o = 32'h00000000 /* 0x11b8 */;
                1135: data_o = 32'h00000000 /* 0x11bc */;
                1136: data_o = 32'h00000000 /* 0x11c0 */;
                1137: data_o = 32'h00000000 /* 0x11c4 */;
                1138: data_o = 32'h00000000 /* 0x11c8 */;
                1139: data_o = 32'h00000000 /* 0x11cc */;
                1140: data_o = 32'h00000000 /* 0x11d0 */;
                1141: data_o = 32'h00000000 /* 0x11d4 */;
                1142: data_o = 32'h00000000 /* 0x11d8 */;
                1143: data_o = 32'h00000000 /* 0x11dc */;
                1144: data_o = 32'h00000000 /* 0x11e0 */;
                1145: data_o = 32'h00000000 /* 0x11e4 */;
                1146: data_o = 32'h00000000 /* 0x11e8 */;
                1147: data_o = 32'h00000000 /* 0x11ec */;
                1148: data_o = 32'h00000000 /* 0x11f0 */;
                1149: data_o = 32'h00000000 /* 0x11f4 */;
                1150: data_o = 32'h00000000 /* 0x11f8 */;
                1151: data_o = 32'h00000000 /* 0x11fc */;
                1152: data_o = 32'h00000000 /* 0x1200 */;
                1153: data_o = 32'h00000000 /* 0x1204 */;
                1154: data_o = 32'h00000000 /* 0x1208 */;
                1155: data_o = 32'h00000000 /* 0x120c */;
                1156: data_o = 32'h00000000 /* 0x1210 */;
                1157: data_o = 32'h00000000 /* 0x1214 */;
                1158: data_o = 32'h00000000 /* 0x1218 */;
                1159: data_o = 32'h00000000 /* 0x121c */;
                1160: data_o = 32'h00000000 /* 0x1220 */;
                1161: data_o = 32'h00000000 /* 0x1224 */;
                1162: data_o = 32'h00000000 /* 0x1228 */;
                1163: data_o = 32'h00000000 /* 0x122c */;
                1164: data_o = 32'h00000000 /* 0x1230 */;
                1165: data_o = 32'h00000000 /* 0x1234 */;
                1166: data_o = 32'h00000000 /* 0x1238 */;
                1167: data_o = 32'h00000000 /* 0x123c */;
                1168: data_o = 32'h00000000 /* 0x1240 */;
                1169: data_o = 32'h00000000 /* 0x1244 */;
                1170: data_o = 32'h00000000 /* 0x1248 */;
                1171: data_o = 32'h00000000 /* 0x124c */;
                1172: data_o = 32'h00000000 /* 0x1250 */;
                1173: data_o = 32'h00000000 /* 0x1254 */;
                1174: data_o = 32'h00000000 /* 0x1258 */;
                1175: data_o = 32'h00000000 /* 0x125c */;
                1176: data_o = 32'h00000000 /* 0x1260 */;
                1177: data_o = 32'h00000000 /* 0x1264 */;
                1178: data_o = 32'h00000000 /* 0x1268 */;
                1179: data_o = 32'h00000000 /* 0x126c */;
                1180: data_o = 32'h00000000 /* 0x1270 */;
                1181: data_o = 32'h00000000 /* 0x1274 */;
                1182: data_o = 32'h00000000 /* 0x1278 */;
                1183: data_o = 32'h00000000 /* 0x127c */;
                1184: data_o = 32'h00000000 /* 0x1280 */;
                1185: data_o = 32'h00000000 /* 0x1284 */;
                1186: data_o = 32'h00000000 /* 0x1288 */;
                1187: data_o = 32'h00000000 /* 0x128c */;
                1188: data_o = 32'h00000000 /* 0x1290 */;
                1189: data_o = 32'h00000000 /* 0x1294 */;
                1190: data_o = 32'h00000000 /* 0x1298 */;
                1191: data_o = 32'h00000000 /* 0x129c */;
                1192: data_o = 32'h00000000 /* 0x12a0 */;
                1193: data_o = 32'h00000000 /* 0x12a4 */;
                1194: data_o = 32'h00000000 /* 0x12a8 */;
                1195: data_o = 32'h00000000 /* 0x12ac */;
                1196: data_o = 32'h00000000 /* 0x12b0 */;
                1197: data_o = 32'h00000000 /* 0x12b4 */;
                1198: data_o = 32'h00000000 /* 0x12b8 */;
                1199: data_o = 32'h00000000 /* 0x12bc */;
                1200: data_o = 32'h00000000 /* 0x12c0 */;
                1201: data_o = 32'h00000000 /* 0x12c4 */;
                1202: data_o = 32'h00000000 /* 0x12c8 */;
                1203: data_o = 32'h00000000 /* 0x12cc */;
                1204: data_o = 32'h00000000 /* 0x12d0 */;
                1205: data_o = 32'h00000000 /* 0x12d4 */;
                1206: data_o = 32'h00000000 /* 0x12d8 */;
                1207: data_o = 32'h00000000 /* 0x12dc */;
                1208: data_o = 32'h00000000 /* 0x12e0 */;
                1209: data_o = 32'h00000000 /* 0x12e4 */;
                1210: data_o = 32'h00000000 /* 0x12e8 */;
                1211: data_o = 32'h00000000 /* 0x12ec */;
                1212: data_o = 32'h00000000 /* 0x12f0 */;
                1213: data_o = 32'h00000000 /* 0x12f4 */;
                1214: data_o = 32'h00000000 /* 0x12f8 */;
                1215: data_o = 32'h00000000 /* 0x12fc */;
                1216: data_o = 32'h00000000 /* 0x1300 */;
                1217: data_o = 32'h00000000 /* 0x1304 */;
                1218: data_o = 32'h00000000 /* 0x1308 */;
                1219: data_o = 32'h00000000 /* 0x130c */;
                1220: data_o = 32'h00000000 /* 0x1310 */;
                1221: data_o = 32'h00000000 /* 0x1314 */;
                1222: data_o = 32'h00000000 /* 0x1318 */;
                1223: data_o = 32'h00000000 /* 0x131c */;
                1224: data_o = 32'h00000000 /* 0x1320 */;
                1225: data_o = 32'h00000000 /* 0x1324 */;
                1226: data_o = 32'h00000000 /* 0x1328 */;
                1227: data_o = 32'h00000000 /* 0x132c */;
                1228: data_o = 32'h00000000 /* 0x1330 */;
                1229: data_o = 32'h00000000 /* 0x1334 */;
                1230: data_o = 32'h00000000 /* 0x1338 */;
                1231: data_o = 32'h00000000 /* 0x133c */;
                1232: data_o = 32'h00000000 /* 0x1340 */;
                1233: data_o = 32'h00000000 /* 0x1344 */;
                1234: data_o = 32'h00000000 /* 0x1348 */;
                1235: data_o = 32'h00000000 /* 0x134c */;
                1236: data_o = 32'h00000000 /* 0x1350 */;
                1237: data_o = 32'h00000000 /* 0x1354 */;
                1238: data_o = 32'h00000000 /* 0x1358 */;
                1239: data_o = 32'h00000000 /* 0x135c */;
                1240: data_o = 32'h00000000 /* 0x1360 */;
                1241: data_o = 32'h00000000 /* 0x1364 */;
                1242: data_o = 32'h00000000 /* 0x1368 */;
                1243: data_o = 32'h00000000 /* 0x136c */;
                1244: data_o = 32'h00000000 /* 0x1370 */;
                1245: data_o = 32'h00000000 /* 0x1374 */;
                1246: data_o = 32'h00000000 /* 0x1378 */;
                1247: data_o = 32'h00000000 /* 0x137c */;
                1248: data_o = 32'h00000000 /* 0x1380 */;
                1249: data_o = 32'h00000000 /* 0x1384 */;
                1250: data_o = 32'h00000000 /* 0x1388 */;
                1251: data_o = 32'h00000000 /* 0x138c */;
                1252: data_o = 32'h00000000 /* 0x1390 */;
                1253: data_o = 32'h00000000 /* 0x1394 */;
                1254: data_o = 32'h00000000 /* 0x1398 */;
                1255: data_o = 32'h00000000 /* 0x139c */;
                1256: data_o = 32'h00000000 /* 0x13a0 */;
                1257: data_o = 32'h00000000 /* 0x13a4 */;
                1258: data_o = 32'h00000000 /* 0x13a8 */;
                1259: data_o = 32'h00000000 /* 0x13ac */;
                1260: data_o = 32'h00000000 /* 0x13b0 */;
                1261: data_o = 32'h00000000 /* 0x13b4 */;
                1262: data_o = 32'h00000000 /* 0x13b8 */;
                1263: data_o = 32'h00000000 /* 0x13bc */;
                1264: data_o = 32'h00000000 /* 0x13c0 */;
                1265: data_o = 32'h00000000 /* 0x13c4 */;
                1266: data_o = 32'h00000000 /* 0x13c8 */;
                1267: data_o = 32'h00000000 /* 0x13cc */;
                1268: data_o = 32'h00000000 /* 0x13d0 */;
                1269: data_o = 32'h00000000 /* 0x13d4 */;
                1270: data_o = 32'h00000000 /* 0x13d8 */;
                1271: data_o = 32'h00000000 /* 0x13dc */;
                1272: data_o = 32'h00000000 /* 0x13e0 */;
                1273: data_o = 32'h00000000 /* 0x13e4 */;
                1274: data_o = 32'h00000000 /* 0x13e8 */;
                1275: data_o = 32'h00000000 /* 0x13ec */;
                1276: data_o = 32'h00000000 /* 0x13f0 */;
                1277: data_o = 32'h00000000 /* 0x13f4 */;
                1278: data_o = 32'h00000000 /* 0x13f8 */;
                1279: data_o = 32'h00000000 /* 0x13fc */;
                1280: data_o = 32'h00000000 /* 0x1400 */;
                1281: data_o = 32'h00000000 /* 0x1404 */;
                1282: data_o = 32'h00000000 /* 0x1408 */;
                1283: data_o = 32'h00000000 /* 0x140c */;
                1284: data_o = 32'h00000000 /* 0x1410 */;
                1285: data_o = 32'h00000000 /* 0x1414 */;
                1286: data_o = 32'h00000000 /* 0x1418 */;
                1287: data_o = 32'h00000000 /* 0x141c */;
                1288: data_o = 32'h00000000 /* 0x1420 */;
                1289: data_o = 32'h00000000 /* 0x1424 */;
                1290: data_o = 32'h00000000 /* 0x1428 */;
                1291: data_o = 32'h00000000 /* 0x142c */;
                1292: data_o = 32'h00000000 /* 0x1430 */;
                1293: data_o = 32'h00000000 /* 0x1434 */;
                1294: data_o = 32'h00000000 /* 0x1438 */;
                1295: data_o = 32'h00000000 /* 0x143c */;
                1296: data_o = 32'h00000000 /* 0x1440 */;
                1297: data_o = 32'h00000000 /* 0x1444 */;
                1298: data_o = 32'h00000000 /* 0x1448 */;
                1299: data_o = 32'h00000000 /* 0x144c */;
                1300: data_o = 32'h00000000 /* 0x1450 */;
                1301: data_o = 32'h00000000 /* 0x1454 */;
                1302: data_o = 32'h00000000 /* 0x1458 */;
                1303: data_o = 32'h00000000 /* 0x145c */;
                1304: data_o = 32'h00000000 /* 0x1460 */;
                1305: data_o = 32'h00000000 /* 0x1464 */;
                1306: data_o = 32'h00000000 /* 0x1468 */;
                1307: data_o = 32'h00000000 /* 0x146c */;
                1308: data_o = 32'h00000000 /* 0x1470 */;
                1309: data_o = 32'h00000000 /* 0x1474 */;
                1310: data_o = 32'h00000000 /* 0x1478 */;
                1311: data_o = 32'h00000000 /* 0x147c */;
                1312: data_o = 32'h00000000 /* 0x1480 */;
                1313: data_o = 32'h00000000 /* 0x1484 */;
                1314: data_o = 32'h00000000 /* 0x1488 */;
                1315: data_o = 32'h00000000 /* 0x148c */;
                1316: data_o = 32'h00000000 /* 0x1490 */;
                1317: data_o = 32'h00000000 /* 0x1494 */;
                1318: data_o = 32'h00000000 /* 0x1498 */;
                1319: data_o = 32'h00000000 /* 0x149c */;
                1320: data_o = 32'h00000000 /* 0x14a0 */;
                1321: data_o = 32'h00000000 /* 0x14a4 */;
                1322: data_o = 32'h00000000 /* 0x14a8 */;
                1323: data_o = 32'h00000000 /* 0x14ac */;
                1324: data_o = 32'h00000000 /* 0x14b0 */;
                1325: data_o = 32'h00000000 /* 0x14b4 */;
                1326: data_o = 32'h00000000 /* 0x14b8 */;
                1327: data_o = 32'h00000000 /* 0x14bc */;
                1328: data_o = 32'h00000000 /* 0x14c0 */;
                1329: data_o = 32'h00000000 /* 0x14c4 */;
                1330: data_o = 32'h00000000 /* 0x14c8 */;
                1331: data_o = 32'h00000000 /* 0x14cc */;
                1332: data_o = 32'h00000000 /* 0x14d0 */;
                1333: data_o = 32'h00000000 /* 0x14d4 */;
                1334: data_o = 32'h00000000 /* 0x14d8 */;
                1335: data_o = 32'h00000000 /* 0x14dc */;
                1336: data_o = 32'h00000000 /* 0x14e0 */;
                1337: data_o = 32'h00000000 /* 0x14e4 */;
                1338: data_o = 32'h00000000 /* 0x14e8 */;
                1339: data_o = 32'h00000000 /* 0x14ec */;
                1340: data_o = 32'h00000000 /* 0x14f0 */;
                1341: data_o = 32'h00000000 /* 0x14f4 */;
                1342: data_o = 32'h00000000 /* 0x14f8 */;
                1343: data_o = 32'h00000000 /* 0x14fc */;
                1344: data_o = 32'h00000000 /* 0x1500 */;
                1345: data_o = 32'h00000000 /* 0x1504 */;
                1346: data_o = 32'h00000000 /* 0x1508 */;
                1347: data_o = 32'h00000000 /* 0x150c */;
                1348: data_o = 32'h00000000 /* 0x1510 */;
                1349: data_o = 32'h00000000 /* 0x1514 */;
                1350: data_o = 32'h00000000 /* 0x1518 */;
                1351: data_o = 32'h00000000 /* 0x151c */;
                1352: data_o = 32'h00000000 /* 0x1520 */;
                1353: data_o = 32'h00000000 /* 0x1524 */;
                1354: data_o = 32'h00000000 /* 0x1528 */;
                1355: data_o = 32'h00000000 /* 0x152c */;
                1356: data_o = 32'h00000000 /* 0x1530 */;
                1357: data_o = 32'h00000000 /* 0x1534 */;
                1358: data_o = 32'h00000000 /* 0x1538 */;
                1359: data_o = 32'h00000000 /* 0x153c */;
                1360: data_o = 32'h00000000 /* 0x1540 */;
                1361: data_o = 32'h00000000 /* 0x1544 */;
                1362: data_o = 32'h00000000 /* 0x1548 */;
                1363: data_o = 32'h00000000 /* 0x154c */;
                1364: data_o = 32'h00000000 /* 0x1550 */;
                1365: data_o = 32'h00000000 /* 0x1554 */;
                1366: data_o = 32'h00000000 /* 0x1558 */;
                1367: data_o = 32'h00000000 /* 0x155c */;
                1368: data_o = 32'h00000000 /* 0x1560 */;
                1369: data_o = 32'h00000000 /* 0x1564 */;
                1370: data_o = 32'h00000000 /* 0x1568 */;
                1371: data_o = 32'h00000000 /* 0x156c */;
                1372: data_o = 32'h00000000 /* 0x1570 */;
                1373: data_o = 32'h00000000 /* 0x1574 */;
                1374: data_o = 32'h00000000 /* 0x1578 */;
                1375: data_o = 32'h00000000 /* 0x157c */;
                1376: data_o = 32'h00000000 /* 0x1580 */;
                1377: data_o = 32'h00000000 /* 0x1584 */;
                1378: data_o = 32'h00000000 /* 0x1588 */;
                1379: data_o = 32'h00000000 /* 0x158c */;
                1380: data_o = 32'h00000000 /* 0x1590 */;
                1381: data_o = 32'h00000000 /* 0x1594 */;
                1382: data_o = 32'h00000000 /* 0x1598 */;
                1383: data_o = 32'h00000000 /* 0x159c */;
                1384: data_o = 32'h00000000 /* 0x15a0 */;
                1385: data_o = 32'h00000000 /* 0x15a4 */;
                1386: data_o = 32'h00000000 /* 0x15a8 */;
                1387: data_o = 32'h00000000 /* 0x15ac */;
                1388: data_o = 32'h00000000 /* 0x15b0 */;
                1389: data_o = 32'h00000000 /* 0x15b4 */;
                1390: data_o = 32'h00000000 /* 0x15b8 */;
                1391: data_o = 32'h00000000 /* 0x15bc */;
                1392: data_o = 32'h00000000 /* 0x15c0 */;
                1393: data_o = 32'h00000000 /* 0x15c4 */;
                1394: data_o = 32'h00000000 /* 0x15c8 */;
                1395: data_o = 32'h00000000 /* 0x15cc */;
                1396: data_o = 32'h00000000 /* 0x15d0 */;
                1397: data_o = 32'h00000000 /* 0x15d4 */;
                1398: data_o = 32'h00000000 /* 0x15d8 */;
                1399: data_o = 32'h00000000 /* 0x15dc */;
                1400: data_o = 32'h00000000 /* 0x15e0 */;
                1401: data_o = 32'h00000000 /* 0x15e4 */;
                1402: data_o = 32'h00000000 /* 0x15e8 */;
                1403: data_o = 32'h00000000 /* 0x15ec */;
                1404: data_o = 32'h00000000 /* 0x15f0 */;
                1405: data_o = 32'h00000000 /* 0x15f4 */;
                1406: data_o = 32'h00000000 /* 0x15f8 */;
                1407: data_o = 32'h00000000 /* 0x15fc */;
                1408: data_o = 32'h00000000 /* 0x1600 */;
                1409: data_o = 32'h00000000 /* 0x1604 */;
                1410: data_o = 32'h00000000 /* 0x1608 */;
                1411: data_o = 32'h00000000 /* 0x160c */;
                1412: data_o = 32'h00000000 /* 0x1610 */;
                1413: data_o = 32'h00000000 /* 0x1614 */;
                1414: data_o = 32'h00000000 /* 0x1618 */;
                1415: data_o = 32'h00000000 /* 0x161c */;
                1416: data_o = 32'h00000000 /* 0x1620 */;
                1417: data_o = 32'h00000000 /* 0x1624 */;
                1418: data_o = 32'h00000000 /* 0x1628 */;
                1419: data_o = 32'h00000000 /* 0x162c */;
                1420: data_o = 32'h00000000 /* 0x1630 */;
                1421: data_o = 32'h00000000 /* 0x1634 */;
                1422: data_o = 32'h00000000 /* 0x1638 */;
                1423: data_o = 32'h00000000 /* 0x163c */;
                1424: data_o = 32'h00000000 /* 0x1640 */;
                1425: data_o = 32'h00000000 /* 0x1644 */;
                1426: data_o = 32'h00000000 /* 0x1648 */;
                1427: data_o = 32'h00000000 /* 0x164c */;
                1428: data_o = 32'h00000000 /* 0x1650 */;
                1429: data_o = 32'h00000000 /* 0x1654 */;
                1430: data_o = 32'h00000000 /* 0x1658 */;
                1431: data_o = 32'h00000000 /* 0x165c */;
                1432: data_o = 32'h00000000 /* 0x1660 */;
                1433: data_o = 32'h00000000 /* 0x1664 */;
                1434: data_o = 32'h00000000 /* 0x1668 */;
                1435: data_o = 32'h00000000 /* 0x166c */;
                1436: data_o = 32'h00000000 /* 0x1670 */;
                1437: data_o = 32'h00000000 /* 0x1674 */;
                1438: data_o = 32'h00000000 /* 0x1678 */;
                1439: data_o = 32'h00000000 /* 0x167c */;
                1440: data_o = 32'h00000000 /* 0x1680 */;
                1441: data_o = 32'h00000000 /* 0x1684 */;
                1442: data_o = 32'h00000000 /* 0x1688 */;
                1443: data_o = 32'h00000000 /* 0x168c */;
                1444: data_o = 32'h00000000 /* 0x1690 */;
                1445: data_o = 32'h00000000 /* 0x1694 */;
                1446: data_o = 32'h00000000 /* 0x1698 */;
                1447: data_o = 32'h00000000 /* 0x169c */;
                1448: data_o = 32'h00000000 /* 0x16a0 */;
                1449: data_o = 32'h00000000 /* 0x16a4 */;
                1450: data_o = 32'h00000000 /* 0x16a8 */;
                1451: data_o = 32'h00000000 /* 0x16ac */;
                1452: data_o = 32'h00000000 /* 0x16b0 */;
                1453: data_o = 32'h00000000 /* 0x16b4 */;
                1454: data_o = 32'h00000000 /* 0x16b8 */;
                1455: data_o = 32'h00000000 /* 0x16bc */;
                1456: data_o = 32'h00000000 /* 0x16c0 */;
                1457: data_o = 32'h00000000 /* 0x16c4 */;
                1458: data_o = 32'h00000000 /* 0x16c8 */;
                1459: data_o = 32'h00000000 /* 0x16cc */;
                1460: data_o = 32'h00000000 /* 0x16d0 */;
                1461: data_o = 32'h00000000 /* 0x16d4 */;
                1462: data_o = 32'h00000000 /* 0x16d8 */;
                1463: data_o = 32'h00000000 /* 0x16dc */;
                1464: data_o = 32'h00000000 /* 0x16e0 */;
                1465: data_o = 32'h00000000 /* 0x16e4 */;
                1466: data_o = 32'h00000000 /* 0x16e8 */;
                1467: data_o = 32'h00000000 /* 0x16ec */;
                1468: data_o = 32'h00000000 /* 0x16f0 */;
                1469: data_o = 32'h00000000 /* 0x16f4 */;
                1470: data_o = 32'h00000000 /* 0x16f8 */;
                1471: data_o = 32'h00000000 /* 0x16fc */;
                1472: data_o = 32'h00000000 /* 0x1700 */;
                1473: data_o = 32'h00000000 /* 0x1704 */;
                1474: data_o = 32'h00000000 /* 0x1708 */;
                1475: data_o = 32'h00000000 /* 0x170c */;
                1476: data_o = 32'h00000000 /* 0x1710 */;
                1477: data_o = 32'h00000000 /* 0x1714 */;
                1478: data_o = 32'h00000000 /* 0x1718 */;
                1479: data_o = 32'h00000000 /* 0x171c */;
                1480: data_o = 32'h00000000 /* 0x1720 */;
                1481: data_o = 32'h00000000 /* 0x1724 */;
                1482: data_o = 32'h00000000 /* 0x1728 */;
                1483: data_o = 32'h00000000 /* 0x172c */;
                1484: data_o = 32'h00000000 /* 0x1730 */;
                1485: data_o = 32'h00000000 /* 0x1734 */;
                1486: data_o = 32'h00000000 /* 0x1738 */;
                1487: data_o = 32'h00000000 /* 0x173c */;
                1488: data_o = 32'h00000000 /* 0x1740 */;
                1489: data_o = 32'h00000000 /* 0x1744 */;
                1490: data_o = 32'h00000000 /* 0x1748 */;
                1491: data_o = 32'h00000000 /* 0x174c */;
                1492: data_o = 32'h00000000 /* 0x1750 */;
                1493: data_o = 32'h00000000 /* 0x1754 */;
                1494: data_o = 32'h00000000 /* 0x1758 */;
                1495: data_o = 32'h00000000 /* 0x175c */;
                1496: data_o = 32'h00000000 /* 0x1760 */;
                1497: data_o = 32'h00000000 /* 0x1764 */;
                1498: data_o = 32'h00000000 /* 0x1768 */;
                1499: data_o = 32'h00000000 /* 0x176c */;
                1500: data_o = 32'h00000000 /* 0x1770 */;
                1501: data_o = 32'h00000000 /* 0x1774 */;
                1502: data_o = 32'h00000000 /* 0x1778 */;
                1503: data_o = 32'h00000000 /* 0x177c */;
                1504: data_o = 32'h00000000 /* 0x1780 */;
                1505: data_o = 32'h00000000 /* 0x1784 */;
                1506: data_o = 32'h00000000 /* 0x1788 */;
                1507: data_o = 32'h00000000 /* 0x178c */;
                1508: data_o = 32'h00000000 /* 0x1790 */;
                1509: data_o = 32'h00000000 /* 0x1794 */;
                1510: data_o = 32'h00000000 /* 0x1798 */;
                1511: data_o = 32'h00000000 /* 0x179c */;
                1512: data_o = 32'h00000000 /* 0x17a0 */;
                1513: data_o = 32'h00000000 /* 0x17a4 */;
                1514: data_o = 32'h00000000 /* 0x17a8 */;
                1515: data_o = 32'h00000000 /* 0x17ac */;
                1516: data_o = 32'h00000000 /* 0x17b0 */;
                1517: data_o = 32'h00000000 /* 0x17b4 */;
                1518: data_o = 32'h00000000 /* 0x17b8 */;
                1519: data_o = 32'h00000000 /* 0x17bc */;
                1520: data_o = 32'h00000000 /* 0x17c0 */;
                1521: data_o = 32'h00000000 /* 0x17c4 */;
                1522: data_o = 32'h00000000 /* 0x17c8 */;
                1523: data_o = 32'h00000000 /* 0x17cc */;
                1524: data_o = 32'h00000000 /* 0x17d0 */;
                1525: data_o = 32'h00000000 /* 0x17d4 */;
                1526: data_o = 32'h00000000 /* 0x17d8 */;
                1527: data_o = 32'h00000000 /* 0x17dc */;
                1528: data_o = 32'h00000000 /* 0x17e0 */;
                1529: data_o = 32'h00000000 /* 0x17e4 */;
                1530: data_o = 32'h00000000 /* 0x17e8 */;
                1531: data_o = 32'h00000000 /* 0x17ec */;
                1532: data_o = 32'h00000000 /* 0x17f0 */;
                1533: data_o = 32'h00000000 /* 0x17f4 */;
                1534: data_o = 32'h00000000 /* 0x17f8 */;
                1535: data_o = 32'h00000000 /* 0x17fc */;
                1536: data_o = 32'h00000000 /* 0x1800 */;
                1537: data_o = 32'h00000000 /* 0x1804 */;
                1538: data_o = 32'h00000000 /* 0x1808 */;
                1539: data_o = 32'h00000000 /* 0x180c */;
                1540: data_o = 32'h00000000 /* 0x1810 */;
                1541: data_o = 32'h00000000 /* 0x1814 */;
                1542: data_o = 32'h00000000 /* 0x1818 */;
                1543: data_o = 32'h00000000 /* 0x181c */;
                1544: data_o = 32'h00000000 /* 0x1820 */;
                1545: data_o = 32'h00000000 /* 0x1824 */;
                1546: data_o = 32'h00000000 /* 0x1828 */;
                1547: data_o = 32'h00000000 /* 0x182c */;
                1548: data_o = 32'h00000000 /* 0x1830 */;
                1549: data_o = 32'h00000000 /* 0x1834 */;
                1550: data_o = 32'h00000000 /* 0x1838 */;
                1551: data_o = 32'h00000000 /* 0x183c */;
                1552: data_o = 32'h00000000 /* 0x1840 */;
                1553: data_o = 32'h00000000 /* 0x1844 */;
                1554: data_o = 32'h00000000 /* 0x1848 */;
                1555: data_o = 32'h00000000 /* 0x184c */;
                1556: data_o = 32'h00000000 /* 0x1850 */;
                1557: data_o = 32'h00000000 /* 0x1854 */;
                1558: data_o = 32'h00000000 /* 0x1858 */;
                1559: data_o = 32'h00000000 /* 0x185c */;
                1560: data_o = 32'h00000000 /* 0x1860 */;
                1561: data_o = 32'h00000000 /* 0x1864 */;
                1562: data_o = 32'h00000000 /* 0x1868 */;
                1563: data_o = 32'h00000000 /* 0x186c */;
                1564: data_o = 32'h00000000 /* 0x1870 */;
                1565: data_o = 32'h00000000 /* 0x1874 */;
                1566: data_o = 32'h00000000 /* 0x1878 */;
                1567: data_o = 32'h00000000 /* 0x187c */;
                1568: data_o = 32'h00000000 /* 0x1880 */;
                1569: data_o = 32'h00000000 /* 0x1884 */;
                1570: data_o = 32'h00000000 /* 0x1888 */;
                1571: data_o = 32'h00000000 /* 0x188c */;
                1572: data_o = 32'h00000000 /* 0x1890 */;
                1573: data_o = 32'h00000000 /* 0x1894 */;
                1574: data_o = 32'h00000000 /* 0x1898 */;
                1575: data_o = 32'h00000000 /* 0x189c */;
                1576: data_o = 32'h00000000 /* 0x18a0 */;
                1577: data_o = 32'h00000000 /* 0x18a4 */;
                1578: data_o = 32'h00000000 /* 0x18a8 */;
                1579: data_o = 32'h00000000 /* 0x18ac */;
                1580: data_o = 32'h00000000 /* 0x18b0 */;
                1581: data_o = 32'h00000000 /* 0x18b4 */;
                1582: data_o = 32'h00000000 /* 0x18b8 */;
                1583: data_o = 32'h00000000 /* 0x18bc */;
                1584: data_o = 32'h00000000 /* 0x18c0 */;
                1585: data_o = 32'h00000000 /* 0x18c4 */;
                1586: data_o = 32'h00000000 /* 0x18c8 */;
                1587: data_o = 32'h00000000 /* 0x18cc */;
                1588: data_o = 32'h00000000 /* 0x18d0 */;
                1589: data_o = 32'h00000000 /* 0x18d4 */;
                1590: data_o = 32'h00000000 /* 0x18d8 */;
                1591: data_o = 32'h00000000 /* 0x18dc */;
                1592: data_o = 32'h00000000 /* 0x18e0 */;
                1593: data_o = 32'h00000000 /* 0x18e4 */;
                1594: data_o = 32'h00000000 /* 0x18e8 */;
                1595: data_o = 32'h00000000 /* 0x18ec */;
                1596: data_o = 32'h00000000 /* 0x18f0 */;
                1597: data_o = 32'h00000000 /* 0x18f4 */;
                1598: data_o = 32'h00000000 /* 0x18f8 */;
                1599: data_o = 32'h00000000 /* 0x18fc */;
                1600: data_o = 32'h00000000 /* 0x1900 */;
                1601: data_o = 32'h00000000 /* 0x1904 */;
                1602: data_o = 32'h00000000 /* 0x1908 */;
                1603: data_o = 32'h00000000 /* 0x190c */;
                1604: data_o = 32'h00000000 /* 0x1910 */;
                1605: data_o = 32'h00000000 /* 0x1914 */;
                1606: data_o = 32'h00000000 /* 0x1918 */;
                1607: data_o = 32'h00000000 /* 0x191c */;
                1608: data_o = 32'h00000000 /* 0x1920 */;
                1609: data_o = 32'h00000000 /* 0x1924 */;
                1610: data_o = 32'h00000000 /* 0x1928 */;
                1611: data_o = 32'h00000000 /* 0x192c */;
                1612: data_o = 32'h00000000 /* 0x1930 */;
                1613: data_o = 32'h00000000 /* 0x1934 */;
                1614: data_o = 32'h00000000 /* 0x1938 */;
                1615: data_o = 32'h00000000 /* 0x193c */;
                1616: data_o = 32'h00000000 /* 0x1940 */;
                1617: data_o = 32'h00000000 /* 0x1944 */;
                1618: data_o = 32'h00000000 /* 0x1948 */;
                1619: data_o = 32'h00000000 /* 0x194c */;
                1620: data_o = 32'h00000000 /* 0x1950 */;
                1621: data_o = 32'h00000000 /* 0x1954 */;
                1622: data_o = 32'h00000000 /* 0x1958 */;
                1623: data_o = 32'h00000000 /* 0x195c */;
                1624: data_o = 32'h00000000 /* 0x1960 */;
                1625: data_o = 32'h00000000 /* 0x1964 */;
                1626: data_o = 32'h00000000 /* 0x1968 */;
                1627: data_o = 32'h00000000 /* 0x196c */;
                1628: data_o = 32'h00000000 /* 0x1970 */;
                1629: data_o = 32'h00000000 /* 0x1974 */;
                1630: data_o = 32'h00000000 /* 0x1978 */;
                1631: data_o = 32'h00000000 /* 0x197c */;
                1632: data_o = 32'h00000000 /* 0x1980 */;
                1633: data_o = 32'h00000000 /* 0x1984 */;
                1634: data_o = 32'h00000000 /* 0x1988 */;
                1635: data_o = 32'h00000000 /* 0x198c */;
                1636: data_o = 32'h00000000 /* 0x1990 */;
                1637: data_o = 32'h00000000 /* 0x1994 */;
                1638: data_o = 32'h00000000 /* 0x1998 */;
                1639: data_o = 32'h00000000 /* 0x199c */;
                1640: data_o = 32'h00000000 /* 0x19a0 */;
                1641: data_o = 32'h00000000 /* 0x19a4 */;
                1642: data_o = 32'h00000000 /* 0x19a8 */;
                1643: data_o = 32'h00000000 /* 0x19ac */;
                1644: data_o = 32'h00000000 /* 0x19b0 */;
                1645: data_o = 32'h00000000 /* 0x19b4 */;
                1646: data_o = 32'h00000000 /* 0x19b8 */;
                1647: data_o = 32'h00000000 /* 0x19bc */;
                1648: data_o = 32'h00000000 /* 0x19c0 */;
                1649: data_o = 32'h00000000 /* 0x19c4 */;
                1650: data_o = 32'h00000000 /* 0x19c8 */;
                1651: data_o = 32'h00000000 /* 0x19cc */;
                1652: data_o = 32'h00000000 /* 0x19d0 */;
                1653: data_o = 32'h00000000 /* 0x19d4 */;
                1654: data_o = 32'h00000000 /* 0x19d8 */;
                1655: data_o = 32'h00000000 /* 0x19dc */;
                1656: data_o = 32'h00000000 /* 0x19e0 */;
                1657: data_o = 32'h00000000 /* 0x19e4 */;
                1658: data_o = 32'h00000000 /* 0x19e8 */;
                1659: data_o = 32'h00000000 /* 0x19ec */;
                1660: data_o = 32'h00000000 /* 0x19f0 */;
                1661: data_o = 32'h00000000 /* 0x19f4 */;
                1662: data_o = 32'h00000000 /* 0x19f8 */;
                1663: data_o = 32'h00000000 /* 0x19fc */;
                1664: data_o = 32'h00000000 /* 0x1a00 */;
                1665: data_o = 32'h00000000 /* 0x1a04 */;
                1666: data_o = 32'h00000000 /* 0x1a08 */;
                1667: data_o = 32'h00000000 /* 0x1a0c */;
                1668: data_o = 32'h00000000 /* 0x1a10 */;
                1669: data_o = 32'h00000000 /* 0x1a14 */;
                1670: data_o = 32'h00000000 /* 0x1a18 */;
                1671: data_o = 32'h00000000 /* 0x1a1c */;
                1672: data_o = 32'h00000000 /* 0x1a20 */;
                1673: data_o = 32'h00000000 /* 0x1a24 */;
                1674: data_o = 32'h00000000 /* 0x1a28 */;
                1675: data_o = 32'h00000000 /* 0x1a2c */;
                1676: data_o = 32'h00000000 /* 0x1a30 */;
                1677: data_o = 32'h00000000 /* 0x1a34 */;
                1678: data_o = 32'h00000000 /* 0x1a38 */;
                1679: data_o = 32'h00000000 /* 0x1a3c */;
                1680: data_o = 32'h00000000 /* 0x1a40 */;
                1681: data_o = 32'h00000000 /* 0x1a44 */;
                1682: data_o = 32'h00000000 /* 0x1a48 */;
                1683: data_o = 32'h00000000 /* 0x1a4c */;
                1684: data_o = 32'h00000000 /* 0x1a50 */;
                1685: data_o = 32'h00000000 /* 0x1a54 */;
                1686: data_o = 32'h00000000 /* 0x1a58 */;
                1687: data_o = 32'h00000000 /* 0x1a5c */;
                1688: data_o = 32'h00000000 /* 0x1a60 */;
                1689: data_o = 32'h00000000 /* 0x1a64 */;
                1690: data_o = 32'h00000000 /* 0x1a68 */;
                1691: data_o = 32'h00000000 /* 0x1a6c */;
                1692: data_o = 32'h00000000 /* 0x1a70 */;
                1693: data_o = 32'h00000000 /* 0x1a74 */;
                1694: data_o = 32'h00000000 /* 0x1a78 */;
                1695: data_o = 32'h00000000 /* 0x1a7c */;
                1696: data_o = 32'h00000000 /* 0x1a80 */;
                1697: data_o = 32'h00000000 /* 0x1a84 */;
                1698: data_o = 32'h00000000 /* 0x1a88 */;
                1699: data_o = 32'h00000000 /* 0x1a8c */;
                1700: data_o = 32'h00000000 /* 0x1a90 */;
                1701: data_o = 32'h00000000 /* 0x1a94 */;
                1702: data_o = 32'h00000000 /* 0x1a98 */;
                1703: data_o = 32'h00000000 /* 0x1a9c */;
                1704: data_o = 32'h00000000 /* 0x1aa0 */;
                1705: data_o = 32'h00000000 /* 0x1aa4 */;
                1706: data_o = 32'h00000000 /* 0x1aa8 */;
                1707: data_o = 32'h00000000 /* 0x1aac */;
                1708: data_o = 32'h00000000 /* 0x1ab0 */;
                1709: data_o = 32'h00000000 /* 0x1ab4 */;
                1710: data_o = 32'h00000000 /* 0x1ab8 */;
                1711: data_o = 32'h00000000 /* 0x1abc */;
                1712: data_o = 32'h00000000 /* 0x1ac0 */;
                1713: data_o = 32'h00000000 /* 0x1ac4 */;
                1714: data_o = 32'h00000000 /* 0x1ac8 */;
                1715: data_o = 32'h00000000 /* 0x1acc */;
                1716: data_o = 32'h00000000 /* 0x1ad0 */;
                1717: data_o = 32'h00000000 /* 0x1ad4 */;
                1718: data_o = 32'h00000000 /* 0x1ad8 */;
                1719: data_o = 32'h00000000 /* 0x1adc */;
                1720: data_o = 32'h00000000 /* 0x1ae0 */;
                1721: data_o = 32'h00000000 /* 0x1ae4 */;
                1722: data_o = 32'h00000000 /* 0x1ae8 */;
                1723: data_o = 32'h00000000 /* 0x1aec */;
                1724: data_o = 32'h00000000 /* 0x1af0 */;
                1725: data_o = 32'h00000000 /* 0x1af4 */;
                1726: data_o = 32'h00000000 /* 0x1af8 */;
                1727: data_o = 32'h00000000 /* 0x1afc */;
                1728: data_o = 32'h00000000 /* 0x1b00 */;
                1729: data_o = 32'h00000000 /* 0x1b04 */;
                1730: data_o = 32'h00000000 /* 0x1b08 */;
                1731: data_o = 32'h00000000 /* 0x1b0c */;
                1732: data_o = 32'h00000000 /* 0x1b10 */;
                1733: data_o = 32'h00000000 /* 0x1b14 */;
                1734: data_o = 32'h00000000 /* 0x1b18 */;
                1735: data_o = 32'h00000000 /* 0x1b1c */;
                1736: data_o = 32'h00000000 /* 0x1b20 */;
                1737: data_o = 32'h00000000 /* 0x1b24 */;
                1738: data_o = 32'h00000000 /* 0x1b28 */;
                1739: data_o = 32'h00000000 /* 0x1b2c */;
                1740: data_o = 32'h00000000 /* 0x1b30 */;
                1741: data_o = 32'h00000000 /* 0x1b34 */;
                1742: data_o = 32'h00000000 /* 0x1b38 */;
                1743: data_o = 32'h00000000 /* 0x1b3c */;
                1744: data_o = 32'h00000000 /* 0x1b40 */;
                1745: data_o = 32'h00000000 /* 0x1b44 */;
                1746: data_o = 32'h00000000 /* 0x1b48 */;
                1747: data_o = 32'h00000000 /* 0x1b4c */;
                1748: data_o = 32'h00000000 /* 0x1b50 */;
                1749: data_o = 32'h00000000 /* 0x1b54 */;
                1750: data_o = 32'h00000000 /* 0x1b58 */;
                1751: data_o = 32'h00000000 /* 0x1b5c */;
                1752: data_o = 32'h00000000 /* 0x1b60 */;
                1753: data_o = 32'h00000000 /* 0x1b64 */;
                1754: data_o = 32'h00000000 /* 0x1b68 */;
                1755: data_o = 32'h00000000 /* 0x1b6c */;
                1756: data_o = 32'h00000000 /* 0x1b70 */;
                1757: data_o = 32'h00000000 /* 0x1b74 */;
                1758: data_o = 32'h00000000 /* 0x1b78 */;
                1759: data_o = 32'h00000000 /* 0x1b7c */;
                1760: data_o = 32'h00000000 /* 0x1b80 */;
                1761: data_o = 32'h00000000 /* 0x1b84 */;
                1762: data_o = 32'h00000000 /* 0x1b88 */;
                1763: data_o = 32'h00000000 /* 0x1b8c */;
                1764: data_o = 32'h00000000 /* 0x1b90 */;
                1765: data_o = 32'h00000000 /* 0x1b94 */;
                1766: data_o = 32'h00000000 /* 0x1b98 */;
                1767: data_o = 32'h00000000 /* 0x1b9c */;
                1768: data_o = 32'h00000000 /* 0x1ba0 */;
                1769: data_o = 32'h00000000 /* 0x1ba4 */;
                1770: data_o = 32'h00000000 /* 0x1ba8 */;
                1771: data_o = 32'h00000000 /* 0x1bac */;
                1772: data_o = 32'h00000000 /* 0x1bb0 */;
                1773: data_o = 32'h00000000 /* 0x1bb4 */;
                1774: data_o = 32'h00000000 /* 0x1bb8 */;
                1775: data_o = 32'h00000000 /* 0x1bbc */;
                1776: data_o = 32'h00000000 /* 0x1bc0 */;
                1777: data_o = 32'h00000000 /* 0x1bc4 */;
                1778: data_o = 32'h00000000 /* 0x1bc8 */;
                1779: data_o = 32'h00000000 /* 0x1bcc */;
                1780: data_o = 32'h00000000 /* 0x1bd0 */;
                1781: data_o = 32'h00000000 /* 0x1bd4 */;
                1782: data_o = 32'h00000000 /* 0x1bd8 */;
                1783: data_o = 32'h00000000 /* 0x1bdc */;
                1784: data_o = 32'h00000000 /* 0x1be0 */;
                1785: data_o = 32'h00000000 /* 0x1be4 */;
                1786: data_o = 32'h00000000 /* 0x1be8 */;
                1787: data_o = 32'h00000000 /* 0x1bec */;
                1788: data_o = 32'h00000000 /* 0x1bf0 */;
                1789: data_o = 32'h00000000 /* 0x1bf4 */;
                1790: data_o = 32'h00000000 /* 0x1bf8 */;
                1791: data_o = 32'h00000000 /* 0x1bfc */;
                1792: data_o = 32'h00000000 /* 0x1c00 */;
                1793: data_o = 32'h00000000 /* 0x1c04 */;
                1794: data_o = 32'h00000000 /* 0x1c08 */;
                1795: data_o = 32'h00000000 /* 0x1c0c */;
                1796: data_o = 32'h00000000 /* 0x1c10 */;
                1797: data_o = 32'h00000000 /* 0x1c14 */;
                1798: data_o = 32'h00000000 /* 0x1c18 */;
                1799: data_o = 32'h00000000 /* 0x1c1c */;
                1800: data_o = 32'h00000000 /* 0x1c20 */;
                1801: data_o = 32'h00000000 /* 0x1c24 */;
                1802: data_o = 32'h00000000 /* 0x1c28 */;
                1803: data_o = 32'h00000000 /* 0x1c2c */;
                1804: data_o = 32'h00000000 /* 0x1c30 */;
                1805: data_o = 32'h00000000 /* 0x1c34 */;
                1806: data_o = 32'h00000000 /* 0x1c38 */;
                1807: data_o = 32'h00000000 /* 0x1c3c */;
                1808: data_o = 32'h00000000 /* 0x1c40 */;
                1809: data_o = 32'h00000000 /* 0x1c44 */;
                1810: data_o = 32'h00000000 /* 0x1c48 */;
                1811: data_o = 32'h00000000 /* 0x1c4c */;
                1812: data_o = 32'h00000000 /* 0x1c50 */;
                1813: data_o = 32'h00000000 /* 0x1c54 */;
                1814: data_o = 32'h00000000 /* 0x1c58 */;
                1815: data_o = 32'h00000000 /* 0x1c5c */;
                1816: data_o = 32'h00000000 /* 0x1c60 */;
                1817: data_o = 32'h00000000 /* 0x1c64 */;
                1818: data_o = 32'h00000000 /* 0x1c68 */;
                1819: data_o = 32'h00000000 /* 0x1c6c */;
                1820: data_o = 32'h00000000 /* 0x1c70 */;
                1821: data_o = 32'h00000000 /* 0x1c74 */;
                1822: data_o = 32'h00000000 /* 0x1c78 */;
                1823: data_o = 32'h00000000 /* 0x1c7c */;
                1824: data_o = 32'h00000000 /* 0x1c80 */;
                1825: data_o = 32'h00000000 /* 0x1c84 */;
                1826: data_o = 32'h00000000 /* 0x1c88 */;
                1827: data_o = 32'h00000000 /* 0x1c8c */;
                1828: data_o = 32'h00000000 /* 0x1c90 */;
                1829: data_o = 32'h00000000 /* 0x1c94 */;
                1830: data_o = 32'h00000000 /* 0x1c98 */;
                1831: data_o = 32'h00000000 /* 0x1c9c */;
                1832: data_o = 32'h00000000 /* 0x1ca0 */;
                1833: data_o = 32'h00000000 /* 0x1ca4 */;
                1834: data_o = 32'h00000000 /* 0x1ca8 */;
                1835: data_o = 32'h00000000 /* 0x1cac */;
                1836: data_o = 32'h00000000 /* 0x1cb0 */;
                1837: data_o = 32'h00000000 /* 0x1cb4 */;
                1838: data_o = 32'h00000000 /* 0x1cb8 */;
                1839: data_o = 32'h00000000 /* 0x1cbc */;
                1840: data_o = 32'h00000000 /* 0x1cc0 */;
                1841: data_o = 32'h00000000 /* 0x1cc4 */;
                1842: data_o = 32'h00000000 /* 0x1cc8 */;
                1843: data_o = 32'h00000000 /* 0x1ccc */;
                1844: data_o = 32'h00000000 /* 0x1cd0 */;
                1845: data_o = 32'h00000000 /* 0x1cd4 */;
                1846: data_o = 32'h00000000 /* 0x1cd8 */;
                1847: data_o = 32'h00000000 /* 0x1cdc */;
                1848: data_o = 32'h00000000 /* 0x1ce0 */;
                1849: data_o = 32'h00000000 /* 0x1ce4 */;
                1850: data_o = 32'h00000000 /* 0x1ce8 */;
                1851: data_o = 32'h00000000 /* 0x1cec */;
                1852: data_o = 32'h00000000 /* 0x1cf0 */;
                1853: data_o = 32'h00000000 /* 0x1cf4 */;
                1854: data_o = 32'h00000000 /* 0x1cf8 */;
                1855: data_o = 32'h00000000 /* 0x1cfc */;
                1856: data_o = 32'h00000000 /* 0x1d00 */;
                1857: data_o = 32'h00000000 /* 0x1d04 */;
                1858: data_o = 32'h00000000 /* 0x1d08 */;
                1859: data_o = 32'h00000000 /* 0x1d0c */;
                1860: data_o = 32'h00000000 /* 0x1d10 */;
                1861: data_o = 32'h00000000 /* 0x1d14 */;
                1862: data_o = 32'h00000000 /* 0x1d18 */;
                1863: data_o = 32'h00000000 /* 0x1d1c */;
                1864: data_o = 32'h00000000 /* 0x1d20 */;
                1865: data_o = 32'h00000000 /* 0x1d24 */;
                1866: data_o = 32'h00000000 /* 0x1d28 */;
                1867: data_o = 32'h00000000 /* 0x1d2c */;
                1868: data_o = 32'h00000000 /* 0x1d30 */;
                1869: data_o = 32'h00000000 /* 0x1d34 */;
                1870: data_o = 32'h00000000 /* 0x1d38 */;
                1871: data_o = 32'h00000000 /* 0x1d3c */;
                1872: data_o = 32'h00000000 /* 0x1d40 */;
                1873: data_o = 32'h00000000 /* 0x1d44 */;
                1874: data_o = 32'h00000000 /* 0x1d48 */;
                1875: data_o = 32'h00000000 /* 0x1d4c */;
                1876: data_o = 32'h00000000 /* 0x1d50 */;
                1877: data_o = 32'h00000000 /* 0x1d54 */;
                1878: data_o = 32'h00000000 /* 0x1d58 */;
                1879: data_o = 32'h00000000 /* 0x1d5c */;
                1880: data_o = 32'h00000000 /* 0x1d60 */;
                1881: data_o = 32'h00000000 /* 0x1d64 */;
                1882: data_o = 32'h00000000 /* 0x1d68 */;
                1883: data_o = 32'h00000000 /* 0x1d6c */;
                1884: data_o = 32'h00000000 /* 0x1d70 */;
                1885: data_o = 32'h00000000 /* 0x1d74 */;
                1886: data_o = 32'h00000000 /* 0x1d78 */;
                1887: data_o = 32'h00000000 /* 0x1d7c */;
                1888: data_o = 32'h00000000 /* 0x1d80 */;
                1889: data_o = 32'h00000000 /* 0x1d84 */;
                1890: data_o = 32'h00000000 /* 0x1d88 */;
                1891: data_o = 32'h00000000 /* 0x1d8c */;
                1892: data_o = 32'h00000000 /* 0x1d90 */;
                1893: data_o = 32'h00000000 /* 0x1d94 */;
                1894: data_o = 32'h00000000 /* 0x1d98 */;
                1895: data_o = 32'h00000000 /* 0x1d9c */;
                1896: data_o = 32'h00000000 /* 0x1da0 */;
                1897: data_o = 32'h00000000 /* 0x1da4 */;
                1898: data_o = 32'h00000000 /* 0x1da8 */;
                1899: data_o = 32'h00000000 /* 0x1dac */;
                1900: data_o = 32'h00000000 /* 0x1db0 */;
                1901: data_o = 32'h00000000 /* 0x1db4 */;
                1902: data_o = 32'h00000000 /* 0x1db8 */;
                1903: data_o = 32'h00000000 /* 0x1dbc */;
                1904: data_o = 32'h00000000 /* 0x1dc0 */;
                1905: data_o = 32'h00000000 /* 0x1dc4 */;
                1906: data_o = 32'h00000000 /* 0x1dc8 */;
                1907: data_o = 32'h00000000 /* 0x1dcc */;
                1908: data_o = 32'h00000000 /* 0x1dd0 */;
                1909: data_o = 32'h00000000 /* 0x1dd4 */;
                1910: data_o = 32'h00000000 /* 0x1dd8 */;
                1911: data_o = 32'h00000000 /* 0x1ddc */;
                1912: data_o = 32'h00000000 /* 0x1de0 */;
                1913: data_o = 32'h00000000 /* 0x1de4 */;
                1914: data_o = 32'h00000000 /* 0x1de8 */;
                1915: data_o = 32'h00000000 /* 0x1dec */;
                1916: data_o = 32'h00000000 /* 0x1df0 */;
                1917: data_o = 32'h00000000 /* 0x1df4 */;
                1918: data_o = 32'h00000000 /* 0x1df8 */;
                1919: data_o = 32'h00000000 /* 0x1dfc */;
                1920: data_o = 32'h00000000 /* 0x1e00 */;
                1921: data_o = 32'h00000000 /* 0x1e04 */;
                1922: data_o = 32'h00000000 /* 0x1e08 */;
                1923: data_o = 32'h00000000 /* 0x1e0c */;
                1924: data_o = 32'h00000000 /* 0x1e10 */;
                1925: data_o = 32'h00000000 /* 0x1e14 */;
                1926: data_o = 32'h00000000 /* 0x1e18 */;
                1927: data_o = 32'h00000000 /* 0x1e1c */;
                1928: data_o = 32'h00000000 /* 0x1e20 */;
                1929: data_o = 32'h00000000 /* 0x1e24 */;
                1930: data_o = 32'h00000000 /* 0x1e28 */;
                1931: data_o = 32'h00000000 /* 0x1e2c */;
                1932: data_o = 32'h00000000 /* 0x1e30 */;
                1933: data_o = 32'h00000000 /* 0x1e34 */;
                1934: data_o = 32'h00000000 /* 0x1e38 */;
                1935: data_o = 32'h00000000 /* 0x1e3c */;
                1936: data_o = 32'h00000000 /* 0x1e40 */;
                1937: data_o = 32'h00000000 /* 0x1e44 */;
                1938: data_o = 32'h00000000 /* 0x1e48 */;
                1939: data_o = 32'h00000000 /* 0x1e4c */;
                1940: data_o = 32'h00000000 /* 0x1e50 */;
                1941: data_o = 32'h00000000 /* 0x1e54 */;
                1942: data_o = 32'h00000000 /* 0x1e58 */;
                1943: data_o = 32'h00000000 /* 0x1e5c */;
                1944: data_o = 32'h00000000 /* 0x1e60 */;
                1945: data_o = 32'h00000000 /* 0x1e64 */;
                1946: data_o = 32'h00000000 /* 0x1e68 */;
                1947: data_o = 32'h00000000 /* 0x1e6c */;
                1948: data_o = 32'h00000000 /* 0x1e70 */;
                1949: data_o = 32'h00000000 /* 0x1e74 */;
                1950: data_o = 32'h00000000 /* 0x1e78 */;
                1951: data_o = 32'h00000000 /* 0x1e7c */;
                1952: data_o = 32'h00000000 /* 0x1e80 */;
                1953: data_o = 32'h00000000 /* 0x1e84 */;
                1954: data_o = 32'h00000000 /* 0x1e88 */;
                1955: data_o = 32'h00000000 /* 0x1e8c */;
                1956: data_o = 32'h00000000 /* 0x1e90 */;
                1957: data_o = 32'h00000000 /* 0x1e94 */;
                1958: data_o = 32'h00000000 /* 0x1e98 */;
                1959: data_o = 32'h00000000 /* 0x1e9c */;
                1960: data_o = 32'h00000000 /* 0x1ea0 */;
                1961: data_o = 32'h00000000 /* 0x1ea4 */;
                1962: data_o = 32'h00000000 /* 0x1ea8 */;
                1963: data_o = 32'h00000000 /* 0x1eac */;
                1964: data_o = 32'h00000000 /* 0x1eb0 */;
                1965: data_o = 32'h00000000 /* 0x1eb4 */;
                1966: data_o = 32'h00000000 /* 0x1eb8 */;
                1967: data_o = 32'h00000000 /* 0x1ebc */;
                1968: data_o = 32'h00000000 /* 0x1ec0 */;
                1969: data_o = 32'h00000000 /* 0x1ec4 */;
                1970: data_o = 32'h00000000 /* 0x1ec8 */;
                1971: data_o = 32'h00000000 /* 0x1ecc */;
                1972: data_o = 32'h00000000 /* 0x1ed0 */;
                1973: data_o = 32'h00000000 /* 0x1ed4 */;
                1974: data_o = 32'h00000000 /* 0x1ed8 */;
                1975: data_o = 32'h00000000 /* 0x1edc */;
                1976: data_o = 32'h00000000 /* 0x1ee0 */;
                1977: data_o = 32'h00000000 /* 0x1ee4 */;
                1978: data_o = 32'h00000000 /* 0x1ee8 */;
                1979: data_o = 32'h00000000 /* 0x1eec */;
                1980: data_o = 32'h00000000 /* 0x1ef0 */;
                1981: data_o = 32'h00000000 /* 0x1ef4 */;
                1982: data_o = 32'h00000000 /* 0x1ef8 */;
                1983: data_o = 32'h00000000 /* 0x1efc */;
                1984: data_o = 32'h00000000 /* 0x1f00 */;
                1985: data_o = 32'h00000000 /* 0x1f04 */;
                1986: data_o = 32'h00000000 /* 0x1f08 */;
                1987: data_o = 32'h00000000 /* 0x1f0c */;
                1988: data_o = 32'h00000000 /* 0x1f10 */;
                1989: data_o = 32'h00000000 /* 0x1f14 */;
                1990: data_o = 32'h00000000 /* 0x1f18 */;
                1991: data_o = 32'h00000000 /* 0x1f1c */;
                1992: data_o = 32'h00000000 /* 0x1f20 */;
                1993: data_o = 32'h00000000 /* 0x1f24 */;
                1994: data_o = 32'h00000000 /* 0x1f28 */;
                1995: data_o = 32'h00000000 /* 0x1f2c */;
                1996: data_o = 32'h00000000 /* 0x1f30 */;
                1997: data_o = 32'h00000000 /* 0x1f34 */;
                1998: data_o = 32'h00000000 /* 0x1f38 */;
                1999: data_o = 32'h00000000 /* 0x1f3c */;
                2000: data_o = 32'h00000000 /* 0x1f40 */;
                2001: data_o = 32'h00000000 /* 0x1f44 */;
                2002: data_o = 32'h00000000 /* 0x1f48 */;
                2003: data_o = 32'h00000000 /* 0x1f4c */;
                2004: data_o = 32'h00000000 /* 0x1f50 */;
                2005: data_o = 32'h00000000 /* 0x1f54 */;
                2006: data_o = 32'h00000000 /* 0x1f58 */;
                2007: data_o = 32'h00000000 /* 0x1f5c */;
                2008: data_o = 32'h00000000 /* 0x1f60 */;
                2009: data_o = 32'h00000000 /* 0x1f64 */;
                2010: data_o = 32'h00000000 /* 0x1f68 */;
                2011: data_o = 32'h00000000 /* 0x1f6c */;
                2012: data_o = 32'h00000000 /* 0x1f70 */;
                2013: data_o = 32'h00000000 /* 0x1f74 */;
                2014: data_o = 32'h00000000 /* 0x1f78 */;
                2015: data_o = 32'h00000000 /* 0x1f7c */;
                2016: data_o = 32'h00000000 /* 0x1f80 */;
                2017: data_o = 32'h00000000 /* 0x1f84 */;
                2018: data_o = 32'h00000000 /* 0x1f88 */;
                2019: data_o = 32'h00000000 /* 0x1f8c */;
                2020: data_o = 32'h00000000 /* 0x1f90 */;
                2021: data_o = 32'h00000000 /* 0x1f94 */;
                2022: data_o = 32'h00000000 /* 0x1f98 */;
                2023: data_o = 32'h00000000 /* 0x1f9c */;
                2024: data_o = 32'h00000000 /* 0x1fa0 */;
                2025: data_o = 32'h00000000 /* 0x1fa4 */;
                2026: data_o = 32'h00000000 /* 0x1fa8 */;
                2027: data_o = 32'h00000000 /* 0x1fac */;
                2028: data_o = 32'h00000000 /* 0x1fb0 */;
                2029: data_o = 32'h00000000 /* 0x1fb4 */;
                2030: data_o = 32'h00000000 /* 0x1fb8 */;
                2031: data_o = 32'h00000000 /* 0x1fbc */;
                2032: data_o = 32'h00000000 /* 0x1fc0 */;
                2033: data_o = 32'h00000000 /* 0x1fc4 */;
                2034: data_o = 32'h00000000 /* 0x1fc8 */;
                2035: data_o = 32'h00000000 /* 0x1fcc */;
                2036: data_o = 32'h00000000 /* 0x1fd0 */;
                2037: data_o = 32'h00000000 /* 0x1fd4 */;
                2038: data_o = 32'h00000000 /* 0x1fd8 */;
                2039: data_o = 32'h00000000 /* 0x1fdc */;
                2040: data_o = 32'h00000000 /* 0x1fe0 */;
                2041: data_o = 32'h00000000 /* 0x1fe4 */;
                2042: data_o = 32'h00000000 /* 0x1fe8 */;
                2043: data_o = 32'h00000000 /* 0x1fec */;
                2044: data_o = 32'h00000000 /* 0x1ff0 */;
                2045: data_o = 32'h00000000 /* 0x1ff4 */;
                2046: data_o = 32'h00000000 /* 0x1ff8 */;
                2047: data_o = 32'h00000000 /* 0x1ffc */;
                2048: data_o = 32'h00000000 /* 0x2000 */;
                2049: data_o = 32'h00000000 /* 0x2004 */;
                2050: data_o = 32'h00000000 /* 0x2008 */;
                2051: data_o = 32'h00000000 /* 0x200c */;
                2052: data_o = 32'h00000000 /* 0x2010 */;
                2053: data_o = 32'h00000000 /* 0x2014 */;
                2054: data_o = 32'h00000000 /* 0x2018 */;
                2055: data_o = 32'h00000000 /* 0x201c */;
                2056: data_o = 32'h00000000 /* 0x2020 */;
                2057: data_o = 32'h00000000 /* 0x2024 */;
                2058: data_o = 32'h00000000 /* 0x2028 */;
                2059: data_o = 32'h00000000 /* 0x202c */;
                2060: data_o = 32'h00000000 /* 0x2030 */;
                2061: data_o = 32'h00000000 /* 0x2034 */;
                2062: data_o = 32'h00000000 /* 0x2038 */;
                2063: data_o = 32'h00000000 /* 0x203c */;
                2064: data_o = 32'h00000000 /* 0x2040 */;
                2065: data_o = 32'h00000000 /* 0x2044 */;
                2066: data_o = 32'h00000000 /* 0x2048 */;
                2067: data_o = 32'h00000000 /* 0x204c */;
                2068: data_o = 32'h00000000 /* 0x2050 */;
                2069: data_o = 32'h00000000 /* 0x2054 */;
                2070: data_o = 32'h00000000 /* 0x2058 */;
                2071: data_o = 32'h00000000 /* 0x205c */;
                2072: data_o = 32'h00000000 /* 0x2060 */;
                2073: data_o = 32'h00000000 /* 0x2064 */;
                2074: data_o = 32'h00000000 /* 0x2068 */;
                2075: data_o = 32'h00000000 /* 0x206c */;
                2076: data_o = 32'h00000000 /* 0x2070 */;
                2077: data_o = 32'h00000000 /* 0x2074 */;
                2078: data_o = 32'h00000000 /* 0x2078 */;
                2079: data_o = 32'h00000000 /* 0x207c */;
                2080: data_o = 32'h00000000 /* 0x2080 */;
                2081: data_o = 32'h00000000 /* 0x2084 */;
                2082: data_o = 32'h00000000 /* 0x2088 */;
                2083: data_o = 32'h00000000 /* 0x208c */;
                2084: data_o = 32'h00000000 /* 0x2090 */;
                2085: data_o = 32'h00000000 /* 0x2094 */;
                2086: data_o = 32'h00000000 /* 0x2098 */;
                2087: data_o = 32'h00000000 /* 0x209c */;
                2088: data_o = 32'h00000000 /* 0x20a0 */;
                2089: data_o = 32'h00000000 /* 0x20a4 */;
                2090: data_o = 32'h00000000 /* 0x20a8 */;
                2091: data_o = 32'h00000000 /* 0x20ac */;
                2092: data_o = 32'h00000000 /* 0x20b0 */;
                2093: data_o = 32'h00000000 /* 0x20b4 */;
                2094: data_o = 32'h00000000 /* 0x20b8 */;
                2095: data_o = 32'h00000000 /* 0x20bc */;
                2096: data_o = 32'h00000000 /* 0x20c0 */;
                2097: data_o = 32'h00000000 /* 0x20c4 */;
                2098: data_o = 32'h00000000 /* 0x20c8 */;
                2099: data_o = 32'h00000000 /* 0x20cc */;
                2100: data_o = 32'h00000000 /* 0x20d0 */;
                2101: data_o = 32'h00000000 /* 0x20d4 */;
                2102: data_o = 32'h00000000 /* 0x20d8 */;
                2103: data_o = 32'h00000000 /* 0x20dc */;
                2104: data_o = 32'h00000000 /* 0x20e0 */;
                2105: data_o = 32'h00000000 /* 0x20e4 */;
                2106: data_o = 32'h00000000 /* 0x20e8 */;
                2107: data_o = 32'h00000000 /* 0x20ec */;
                2108: data_o = 32'h00000000 /* 0x20f0 */;
                2109: data_o = 32'h00000000 /* 0x20f4 */;
                2110: data_o = 32'h00000000 /* 0x20f8 */;
                2111: data_o = 32'h00000000 /* 0x20fc */;
                2112: data_o = 32'h00000000 /* 0x2100 */;
                2113: data_o = 32'h00000000 /* 0x2104 */;
                2114: data_o = 32'h00000000 /* 0x2108 */;
                2115: data_o = 32'h00000000 /* 0x210c */;
                2116: data_o = 32'h00000000 /* 0x2110 */;
                2117: data_o = 32'h00000000 /* 0x2114 */;
                2118: data_o = 32'h00000000 /* 0x2118 */;
                2119: data_o = 32'h00000000 /* 0x211c */;
                2120: data_o = 32'h00000000 /* 0x2120 */;
                2121: data_o = 32'h00000000 /* 0x2124 */;
                2122: data_o = 32'h00000000 /* 0x2128 */;
                2123: data_o = 32'h00000000 /* 0x212c */;
                2124: data_o = 32'h00000000 /* 0x2130 */;
                2125: data_o = 32'h00000000 /* 0x2134 */;
                2126: data_o = 32'h00000000 /* 0x2138 */;
                2127: data_o = 32'h00000000 /* 0x213c */;
                2128: data_o = 32'h00000000 /* 0x2140 */;
                2129: data_o = 32'h00000000 /* 0x2144 */;
                2130: data_o = 32'h00000000 /* 0x2148 */;
                2131: data_o = 32'h00000000 /* 0x214c */;
                2132: data_o = 32'h00000000 /* 0x2150 */;
                2133: data_o = 32'h00000000 /* 0x2154 */;
                2134: data_o = 32'h00000000 /* 0x2158 */;
                2135: data_o = 32'h00000000 /* 0x215c */;
                2136: data_o = 32'h00000000 /* 0x2160 */;
                2137: data_o = 32'h00000000 /* 0x2164 */;
                2138: data_o = 32'h00000000 /* 0x2168 */;
                2139: data_o = 32'h00000000 /* 0x216c */;
                2140: data_o = 32'h00000000 /* 0x2170 */;
                2141: data_o = 32'h00000000 /* 0x2174 */;
                2142: data_o = 32'h00000000 /* 0x2178 */;
                2143: data_o = 32'h00000000 /* 0x217c */;
                2144: data_o = 32'h00000000 /* 0x2180 */;
                2145: data_o = 32'h00000000 /* 0x2184 */;
                2146: data_o = 32'h00000000 /* 0x2188 */;
                2147: data_o = 32'h00000000 /* 0x218c */;
                2148: data_o = 32'h00000000 /* 0x2190 */;
                2149: data_o = 32'h00000000 /* 0x2194 */;
                2150: data_o = 32'h00000000 /* 0x2198 */;
                2151: data_o = 32'h00000000 /* 0x219c */;
                2152: data_o = 32'h00000000 /* 0x21a0 */;
                2153: data_o = 32'h00000000 /* 0x21a4 */;
                2154: data_o = 32'h00000000 /* 0x21a8 */;
                2155: data_o = 32'h00000000 /* 0x21ac */;
                2156: data_o = 32'h00000000 /* 0x21b0 */;
                2157: data_o = 32'h00000000 /* 0x21b4 */;
                2158: data_o = 32'h00000000 /* 0x21b8 */;
                2159: data_o = 32'h00000000 /* 0x21bc */;
                2160: data_o = 32'h00000000 /* 0x21c0 */;
                2161: data_o = 32'h00000000 /* 0x21c4 */;
                2162: data_o = 32'h00000000 /* 0x21c8 */;
                2163: data_o = 32'h00000000 /* 0x21cc */;
                2164: data_o = 32'h00000000 /* 0x21d0 */;
                2165: data_o = 32'h00000000 /* 0x21d4 */;
                2166: data_o = 32'h00000000 /* 0x21d8 */;
                2167: data_o = 32'h00000000 /* 0x21dc */;
                2168: data_o = 32'h00000000 /* 0x21e0 */;
                2169: data_o = 32'h00000000 /* 0x21e4 */;
                2170: data_o = 32'h00000000 /* 0x21e8 */;
                2171: data_o = 32'h00000000 /* 0x21ec */;
                2172: data_o = 32'h00000000 /* 0x21f0 */;
                2173: data_o = 32'h00000000 /* 0x21f4 */;
                2174: data_o = 32'h00000000 /* 0x21f8 */;
                2175: data_o = 32'h00000000 /* 0x21fc */;
                2176: data_o = 32'h00000000 /* 0x2200 */;
                2177: data_o = 32'h00000000 /* 0x2204 */;
                2178: data_o = 32'h00000000 /* 0x2208 */;
                2179: data_o = 32'h00000000 /* 0x220c */;
                2180: data_o = 32'h00000000 /* 0x2210 */;
                2181: data_o = 32'h00000000 /* 0x2214 */;
                2182: data_o = 32'h00000000 /* 0x2218 */;
                2183: data_o = 32'h00000000 /* 0x221c */;
                2184: data_o = 32'h00000000 /* 0x2220 */;
                2185: data_o = 32'h00000000 /* 0x2224 */;
                2186: data_o = 32'h00000000 /* 0x2228 */;
                2187: data_o = 32'h00000000 /* 0x222c */;
                2188: data_o = 32'h00000000 /* 0x2230 */;
                2189: data_o = 32'h00000000 /* 0x2234 */;
                2190: data_o = 32'h00000000 /* 0x2238 */;
                2191: data_o = 32'h00000000 /* 0x223c */;
                2192: data_o = 32'h00000000 /* 0x2240 */;
                2193: data_o = 32'h00000000 /* 0x2244 */;
                2194: data_o = 32'h00000000 /* 0x2248 */;
                2195: data_o = 32'h00000000 /* 0x224c */;
                2196: data_o = 32'h00000000 /* 0x2250 */;
                2197: data_o = 32'h00000000 /* 0x2254 */;
                2198: data_o = 32'h00000000 /* 0x2258 */;
                2199: data_o = 32'h00000000 /* 0x225c */;
                2200: data_o = 32'h00000000 /* 0x2260 */;
                2201: data_o = 32'h00000000 /* 0x2264 */;
                2202: data_o = 32'h00000000 /* 0x2268 */;
                2203: data_o = 32'h00000000 /* 0x226c */;
                2204: data_o = 32'h00000000 /* 0x2270 */;
                2205: data_o = 32'h00000000 /* 0x2274 */;
                2206: data_o = 32'h00000000 /* 0x2278 */;
                2207: data_o = 32'h00000000 /* 0x227c */;
                2208: data_o = 32'h00000000 /* 0x2280 */;
                2209: data_o = 32'h00000000 /* 0x2284 */;
                2210: data_o = 32'h00000000 /* 0x2288 */;
                2211: data_o = 32'h00000000 /* 0x228c */;
                2212: data_o = 32'h00000000 /* 0x2290 */;
                2213: data_o = 32'h00000000 /* 0x2294 */;
                2214: data_o = 32'h00000000 /* 0x2298 */;
                2215: data_o = 32'h00000000 /* 0x229c */;
                2216: data_o = 32'h00000000 /* 0x22a0 */;
                2217: data_o = 32'h00000000 /* 0x22a4 */;
                2218: data_o = 32'h00000000 /* 0x22a8 */;
                2219: data_o = 32'h00000000 /* 0x22ac */;
                2220: data_o = 32'h00000000 /* 0x22b0 */;
                2221: data_o = 32'h00000000 /* 0x22b4 */;
                2222: data_o = 32'h00000000 /* 0x22b8 */;
                2223: data_o = 32'h00000000 /* 0x22bc */;
                2224: data_o = 32'h00000000 /* 0x22c0 */;
                2225: data_o = 32'h00000000 /* 0x22c4 */;
                2226: data_o = 32'h00000000 /* 0x22c8 */;
                2227: data_o = 32'h00000000 /* 0x22cc */;
                2228: data_o = 32'h00000000 /* 0x22d0 */;
                2229: data_o = 32'h00000000 /* 0x22d4 */;
                2230: data_o = 32'h00000000 /* 0x22d8 */;
                2231: data_o = 32'h00000000 /* 0x22dc */;
                2232: data_o = 32'h00000000 /* 0x22e0 */;
                2233: data_o = 32'h00000000 /* 0x22e4 */;
                2234: data_o = 32'h00000000 /* 0x22e8 */;
                2235: data_o = 32'h00000000 /* 0x22ec */;
                2236: data_o = 32'h00000000 /* 0x22f0 */;
                2237: data_o = 32'h00000000 /* 0x22f4 */;
                2238: data_o = 32'h00000000 /* 0x22f8 */;
                2239: data_o = 32'h00000000 /* 0x22fc */;
                2240: data_o = 32'h00000000 /* 0x2300 */;
                2241: data_o = 32'h00000000 /* 0x2304 */;
                2242: data_o = 32'h00000000 /* 0x2308 */;
                2243: data_o = 32'h00000000 /* 0x230c */;
                2244: data_o = 32'h00000000 /* 0x2310 */;
                2245: data_o = 32'h00000000 /* 0x2314 */;
                2246: data_o = 32'h00000000 /* 0x2318 */;
                2247: data_o = 32'h00000000 /* 0x231c */;
                2248: data_o = 32'h00000000 /* 0x2320 */;
                2249: data_o = 32'h00000000 /* 0x2324 */;
                2250: data_o = 32'h00000000 /* 0x2328 */;
                2251: data_o = 32'h00000000 /* 0x232c */;
                2252: data_o = 32'h00000000 /* 0x2330 */;
                2253: data_o = 32'h00000000 /* 0x2334 */;
                2254: data_o = 32'h00000000 /* 0x2338 */;
                2255: data_o = 32'h00000000 /* 0x233c */;
                2256: data_o = 32'h00000000 /* 0x2340 */;
                2257: data_o = 32'h00000000 /* 0x2344 */;
                2258: data_o = 32'h00000000 /* 0x2348 */;
                2259: data_o = 32'h00000000 /* 0x234c */;
                2260: data_o = 32'h00000000 /* 0x2350 */;
                2261: data_o = 32'h00000000 /* 0x2354 */;
                2262: data_o = 32'h00000000 /* 0x2358 */;
                2263: data_o = 32'h00000000 /* 0x235c */;
                2264: data_o = 32'h00000000 /* 0x2360 */;
                2265: data_o = 32'h00000000 /* 0x2364 */;
                2266: data_o = 32'h00000000 /* 0x2368 */;
                2267: data_o = 32'h00000000 /* 0x236c */;
                2268: data_o = 32'h00000000 /* 0x2370 */;
                2269: data_o = 32'h00000000 /* 0x2374 */;
                2270: data_o = 32'h00000000 /* 0x2378 */;
                2271: data_o = 32'h00000000 /* 0x237c */;
                2272: data_o = 32'h00000000 /* 0x2380 */;
                2273: data_o = 32'h00000000 /* 0x2384 */;
                2274: data_o = 32'h00000000 /* 0x2388 */;
                2275: data_o = 32'h00000000 /* 0x238c */;
                2276: data_o = 32'h00000000 /* 0x2390 */;
                2277: data_o = 32'h00000000 /* 0x2394 */;
                2278: data_o = 32'h00000000 /* 0x2398 */;
                2279: data_o = 32'h00000000 /* 0x239c */;
                2280: data_o = 32'h00000000 /* 0x23a0 */;
                2281: data_o = 32'h00000000 /* 0x23a4 */;
                2282: data_o = 32'h00000000 /* 0x23a8 */;
                2283: data_o = 32'h00000000 /* 0x23ac */;
                2284: data_o = 32'h00000000 /* 0x23b0 */;
                2285: data_o = 32'h00000000 /* 0x23b4 */;
                2286: data_o = 32'h00000000 /* 0x23b8 */;
                2287: data_o = 32'h00000000 /* 0x23bc */;
                2288: data_o = 32'h00000000 /* 0x23c0 */;
                2289: data_o = 32'h00000000 /* 0x23c4 */;
                2290: data_o = 32'h00000000 /* 0x23c8 */;
                2291: data_o = 32'h00000000 /* 0x23cc */;
                2292: data_o = 32'h00000000 /* 0x23d0 */;
                2293: data_o = 32'h00000000 /* 0x23d4 */;
                2294: data_o = 32'h00000000 /* 0x23d8 */;
                2295: data_o = 32'h00000000 /* 0x23dc */;
                2296: data_o = 32'h00000000 /* 0x23e0 */;
                2297: data_o = 32'h00000000 /* 0x23e4 */;
                2298: data_o = 32'h00000000 /* 0x23e8 */;
                2299: data_o = 32'h00000000 /* 0x23ec */;
                2300: data_o = 32'h00000000 /* 0x23f0 */;
                2301: data_o = 32'h00000000 /* 0x23f4 */;
                2302: data_o = 32'h00000000 /* 0x23f8 */;
                2303: data_o = 32'h00000000 /* 0x23fc */;
                2304: data_o = 32'h00000000 /* 0x2400 */;
                2305: data_o = 32'h00000000 /* 0x2404 */;
                2306: data_o = 32'h00000000 /* 0x2408 */;
                2307: data_o = 32'h00000000 /* 0x240c */;
                2308: data_o = 32'h00000000 /* 0x2410 */;
                2309: data_o = 32'h00000000 /* 0x2414 */;
                2310: data_o = 32'h00000000 /* 0x2418 */;
                2311: data_o = 32'h00000000 /* 0x241c */;
                2312: data_o = 32'h00000000 /* 0x2420 */;
                2313: data_o = 32'h00000000 /* 0x2424 */;
                2314: data_o = 32'h00000000 /* 0x2428 */;
                2315: data_o = 32'h00000000 /* 0x242c */;
                2316: data_o = 32'h00000000 /* 0x2430 */;
                2317: data_o = 32'h00000000 /* 0x2434 */;
                2318: data_o = 32'h00000000 /* 0x2438 */;
                2319: data_o = 32'h00000000 /* 0x243c */;
                2320: data_o = 32'h00000000 /* 0x2440 */;
                2321: data_o = 32'h00000000 /* 0x2444 */;
                2322: data_o = 32'h00000000 /* 0x2448 */;
                2323: data_o = 32'h00000000 /* 0x244c */;
                2324: data_o = 32'h00000000 /* 0x2450 */;
                2325: data_o = 32'h00000000 /* 0x2454 */;
                2326: data_o = 32'h00000000 /* 0x2458 */;
                2327: data_o = 32'h00000000 /* 0x245c */;
                2328: data_o = 32'h00000000 /* 0x2460 */;
                2329: data_o = 32'h00000000 /* 0x2464 */;
                2330: data_o = 32'h00000000 /* 0x2468 */;
                2331: data_o = 32'h00000000 /* 0x246c */;
                2332: data_o = 32'h00000000 /* 0x2470 */;
                2333: data_o = 32'h00000000 /* 0x2474 */;
                2334: data_o = 32'h00000000 /* 0x2478 */;
                2335: data_o = 32'h00000000 /* 0x247c */;
                2336: data_o = 32'h00000000 /* 0x2480 */;
                2337: data_o = 32'h00000000 /* 0x2484 */;
                2338: data_o = 32'h00000000 /* 0x2488 */;
                2339: data_o = 32'h00000000 /* 0x248c */;
                2340: data_o = 32'h00000000 /* 0x2490 */;
                2341: data_o = 32'h00000000 /* 0x2494 */;
                2342: data_o = 32'h00000000 /* 0x2498 */;
                2343: data_o = 32'h00000000 /* 0x249c */;
                2344: data_o = 32'h00000000 /* 0x24a0 */;
                2345: data_o = 32'h00000000 /* 0x24a4 */;
                2346: data_o = 32'h00000000 /* 0x24a8 */;
                2347: data_o = 32'h00000000 /* 0x24ac */;
                2348: data_o = 32'h00000000 /* 0x24b0 */;
                2349: data_o = 32'h00000000 /* 0x24b4 */;
                2350: data_o = 32'h00000000 /* 0x24b8 */;
                2351: data_o = 32'h00000000 /* 0x24bc */;
                2352: data_o = 32'h00000000 /* 0x24c0 */;
                2353: data_o = 32'h00000000 /* 0x24c4 */;
                2354: data_o = 32'h00000000 /* 0x24c8 */;
                2355: data_o = 32'h00000000 /* 0x24cc */;
                2356: data_o = 32'h00000000 /* 0x24d0 */;
                2357: data_o = 32'h00000000 /* 0x24d4 */;
                2358: data_o = 32'h00000000 /* 0x24d8 */;
                2359: data_o = 32'h00000000 /* 0x24dc */;
                2360: data_o = 32'h00000000 /* 0x24e0 */;
                2361: data_o = 32'h00000000 /* 0x24e4 */;
                2362: data_o = 32'h00000000 /* 0x24e8 */;
                2363: data_o = 32'h00000000 /* 0x24ec */;
                2364: data_o = 32'h00000000 /* 0x24f0 */;
                2365: data_o = 32'h00000000 /* 0x24f4 */;
                2366: data_o = 32'h00000000 /* 0x24f8 */;
                2367: data_o = 32'h00000000 /* 0x24fc */;
                2368: data_o = 32'h00000000 /* 0x2500 */;
                2369: data_o = 32'h00000000 /* 0x2504 */;
                2370: data_o = 32'h00000000 /* 0x2508 */;
                2371: data_o = 32'h00000000 /* 0x250c */;
                2372: data_o = 32'h00000000 /* 0x2510 */;
                2373: data_o = 32'h00000000 /* 0x2514 */;
                2374: data_o = 32'h00000000 /* 0x2518 */;
                2375: data_o = 32'h00000000 /* 0x251c */;
                2376: data_o = 32'h00000000 /* 0x2520 */;
                2377: data_o = 32'h00000000 /* 0x2524 */;
                2378: data_o = 32'h00000000 /* 0x2528 */;
                2379: data_o = 32'h00000000 /* 0x252c */;
                2380: data_o = 32'h00000000 /* 0x2530 */;
                2381: data_o = 32'h00000000 /* 0x2534 */;
                2382: data_o = 32'h00000000 /* 0x2538 */;
                2383: data_o = 32'h00000000 /* 0x253c */;
                2384: data_o = 32'h00000000 /* 0x2540 */;
                2385: data_o = 32'h00000000 /* 0x2544 */;
                2386: data_o = 32'h00000000 /* 0x2548 */;
                2387: data_o = 32'h00000000 /* 0x254c */;
                2388: data_o = 32'h00000000 /* 0x2550 */;
                2389: data_o = 32'h00000000 /* 0x2554 */;
                2390: data_o = 32'h00000000 /* 0x2558 */;
                2391: data_o = 32'h00000000 /* 0x255c */;
                2392: data_o = 32'h00000000 /* 0x2560 */;
                2393: data_o = 32'h00000000 /* 0x2564 */;
                2394: data_o = 32'h00000000 /* 0x2568 */;
                2395: data_o = 32'h00000000 /* 0x256c */;
                2396: data_o = 32'h00000000 /* 0x2570 */;
                2397: data_o = 32'h00000000 /* 0x2574 */;
                2398: data_o = 32'h00000000 /* 0x2578 */;
                2399: data_o = 32'h00000000 /* 0x257c */;
                2400: data_o = 32'h00000000 /* 0x2580 */;
                2401: data_o = 32'h00000000 /* 0x2584 */;
                2402: data_o = 32'h00000000 /* 0x2588 */;
                2403: data_o = 32'h00000000 /* 0x258c */;
                2404: data_o = 32'h00000000 /* 0x2590 */;
                2405: data_o = 32'h00000000 /* 0x2594 */;
                2406: data_o = 32'h00000000 /* 0x2598 */;
                2407: data_o = 32'h00000000 /* 0x259c */;
                2408: data_o = 32'h00000000 /* 0x25a0 */;
                2409: data_o = 32'h00000000 /* 0x25a4 */;
                2410: data_o = 32'h00000000 /* 0x25a8 */;
                2411: data_o = 32'h00000000 /* 0x25ac */;
                2412: data_o = 32'h00000000 /* 0x25b0 */;
                2413: data_o = 32'h00000000 /* 0x25b4 */;
                2414: data_o = 32'h00000000 /* 0x25b8 */;
                2415: data_o = 32'h00000000 /* 0x25bc */;
                2416: data_o = 32'h00000000 /* 0x25c0 */;
                2417: data_o = 32'h00000000 /* 0x25c4 */;
                2418: data_o = 32'h00000000 /* 0x25c8 */;
                2419: data_o = 32'h00000000 /* 0x25cc */;
                2420: data_o = 32'h00000000 /* 0x25d0 */;
                2421: data_o = 32'h00000000 /* 0x25d4 */;
                2422: data_o = 32'h00000000 /* 0x25d8 */;
                2423: data_o = 32'h00000000 /* 0x25dc */;
                2424: data_o = 32'h00000000 /* 0x25e0 */;
                2425: data_o = 32'h00000000 /* 0x25e4 */;
                2426: data_o = 32'h00000000 /* 0x25e8 */;
                2427: data_o = 32'h00000000 /* 0x25ec */;
                2428: data_o = 32'h00000000 /* 0x25f0 */;
                2429: data_o = 32'h00000000 /* 0x25f4 */;
                2430: data_o = 32'h00000000 /* 0x25f8 */;
                2431: data_o = 32'h00000000 /* 0x25fc */;
                2432: data_o = 32'h00000000 /* 0x2600 */;
                2433: data_o = 32'h00000000 /* 0x2604 */;
                2434: data_o = 32'h00000000 /* 0x2608 */;
                2435: data_o = 32'h00000000 /* 0x260c */;
                2436: data_o = 32'h00000000 /* 0x2610 */;
                2437: data_o = 32'h00000000 /* 0x2614 */;
                2438: data_o = 32'h00000000 /* 0x2618 */;
                2439: data_o = 32'h00000000 /* 0x261c */;
                2440: data_o = 32'h00000000 /* 0x2620 */;
                2441: data_o = 32'h00000000 /* 0x2624 */;
                2442: data_o = 32'h00000000 /* 0x2628 */;
                2443: data_o = 32'h00000000 /* 0x262c */;
                2444: data_o = 32'h00000000 /* 0x2630 */;
                2445: data_o = 32'h00000000 /* 0x2634 */;
                2446: data_o = 32'h00000000 /* 0x2638 */;
                2447: data_o = 32'h00000000 /* 0x263c */;
                2448: data_o = 32'h00000000 /* 0x2640 */;
                2449: data_o = 32'h00000000 /* 0x2644 */;
                2450: data_o = 32'h00000000 /* 0x2648 */;
                2451: data_o = 32'h00000000 /* 0x264c */;
                2452: data_o = 32'h00000000 /* 0x2650 */;
                2453: data_o = 32'h00000000 /* 0x2654 */;
                2454: data_o = 32'h00000000 /* 0x2658 */;
                2455: data_o = 32'h00000000 /* 0x265c */;
                2456: data_o = 32'h00000000 /* 0x2660 */;
                2457: data_o = 32'h00000000 /* 0x2664 */;
                2458: data_o = 32'h00000000 /* 0x2668 */;
                2459: data_o = 32'h00000000 /* 0x266c */;
                2460: data_o = 32'h00000000 /* 0x2670 */;
                2461: data_o = 32'h00000000 /* 0x2674 */;
                2462: data_o = 32'h00000000 /* 0x2678 */;
                2463: data_o = 32'h00000000 /* 0x267c */;
                2464: data_o = 32'h00000000 /* 0x2680 */;
                2465: data_o = 32'h00000000 /* 0x2684 */;
                2466: data_o = 32'h00000000 /* 0x2688 */;
                2467: data_o = 32'h00000000 /* 0x268c */;
                2468: data_o = 32'h00000000 /* 0x2690 */;
                2469: data_o = 32'h00000000 /* 0x2694 */;
                2470: data_o = 32'h00000000 /* 0x2698 */;
                2471: data_o = 32'h00000000 /* 0x269c */;
                2472: data_o = 32'h00000000 /* 0x26a0 */;
                2473: data_o = 32'h00000000 /* 0x26a4 */;
                2474: data_o = 32'h00000000 /* 0x26a8 */;
                2475: data_o = 32'h00000000 /* 0x26ac */;
                2476: data_o = 32'h00000000 /* 0x26b0 */;
                2477: data_o = 32'h00000000 /* 0x26b4 */;
                2478: data_o = 32'h00000000 /* 0x26b8 */;
                2479: data_o = 32'h00000000 /* 0x26bc */;
                2480: data_o = 32'h00000000 /* 0x26c0 */;
                2481: data_o = 32'h00000000 /* 0x26c4 */;
                2482: data_o = 32'h00000000 /* 0x26c8 */;
                2483: data_o = 32'h00000000 /* 0x26cc */;
                2484: data_o = 32'h00000000 /* 0x26d0 */;
                2485: data_o = 32'h00000000 /* 0x26d4 */;
                2486: data_o = 32'h00000000 /* 0x26d8 */;
                2487: data_o = 32'h00000000 /* 0x26dc */;
                2488: data_o = 32'h00000000 /* 0x26e0 */;
                2489: data_o = 32'h00000000 /* 0x26e4 */;
                2490: data_o = 32'h00000000 /* 0x26e8 */;
                2491: data_o = 32'h00000000 /* 0x26ec */;
                2492: data_o = 32'h00000000 /* 0x26f0 */;
                2493: data_o = 32'h00000000 /* 0x26f4 */;
                2494: data_o = 32'h00000000 /* 0x26f8 */;
                2495: data_o = 32'h00000000 /* 0x26fc */;
                2496: data_o = 32'h00000000 /* 0x2700 */;
                2497: data_o = 32'h00000000 /* 0x2704 */;
                2498: data_o = 32'h00000000 /* 0x2708 */;
                2499: data_o = 32'h00000000 /* 0x270c */;
                2500: data_o = 32'h00000000 /* 0x2710 */;
                2501: data_o = 32'h00000000 /* 0x2714 */;
                2502: data_o = 32'h00000000 /* 0x2718 */;
                2503: data_o = 32'h00000000 /* 0x271c */;
                2504: data_o = 32'h00000000 /* 0x2720 */;
                2505: data_o = 32'h00000000 /* 0x2724 */;
                2506: data_o = 32'h00000000 /* 0x2728 */;
                2507: data_o = 32'h00000000 /* 0x272c */;
                2508: data_o = 32'h00000000 /* 0x2730 */;
                2509: data_o = 32'h00000000 /* 0x2734 */;
                2510: data_o = 32'h00000000 /* 0x2738 */;
                2511: data_o = 32'h00000000 /* 0x273c */;
                2512: data_o = 32'h00000000 /* 0x2740 */;
                2513: data_o = 32'h00000000 /* 0x2744 */;
                2514: data_o = 32'h00000000 /* 0x2748 */;
                2515: data_o = 32'h00000000 /* 0x274c */;
                2516: data_o = 32'h00000000 /* 0x2750 */;
                2517: data_o = 32'h00000000 /* 0x2754 */;
                2518: data_o = 32'h00000000 /* 0x2758 */;
                2519: data_o = 32'h00000000 /* 0x275c */;
                2520: data_o = 32'h00000000 /* 0x2760 */;
                2521: data_o = 32'h00000000 /* 0x2764 */;
                2522: data_o = 32'h00000000 /* 0x2768 */;
                2523: data_o = 32'h00000000 /* 0x276c */;
                2524: data_o = 32'h00000000 /* 0x2770 */;
                2525: data_o = 32'h00000000 /* 0x2774 */;
                2526: data_o = 32'h00000000 /* 0x2778 */;
                2527: data_o = 32'h00000000 /* 0x277c */;
                2528: data_o = 32'h00000000 /* 0x2780 */;
                2529: data_o = 32'h00000000 /* 0x2784 */;
                2530: data_o = 32'h00000000 /* 0x2788 */;
                2531: data_o = 32'h00000000 /* 0x278c */;
                2532: data_o = 32'h00000000 /* 0x2790 */;
                2533: data_o = 32'h00000000 /* 0x2794 */;
                2534: data_o = 32'h00000000 /* 0x2798 */;
                2535: data_o = 32'h00000000 /* 0x279c */;
                2536: data_o = 32'h00000000 /* 0x27a0 */;
                2537: data_o = 32'h00000000 /* 0x27a4 */;
                2538: data_o = 32'h00000000 /* 0x27a8 */;
                2539: data_o = 32'h00000000 /* 0x27ac */;
                2540: data_o = 32'h00000000 /* 0x27b0 */;
                2541: data_o = 32'h00000000 /* 0x27b4 */;
                2542: data_o = 32'h00000000 /* 0x27b8 */;
                2543: data_o = 32'h00000000 /* 0x27bc */;
                2544: data_o = 32'h00000000 /* 0x27c0 */;
                2545: data_o = 32'h00000000 /* 0x27c4 */;
                2546: data_o = 32'h00000000 /* 0x27c8 */;
                2547: data_o = 32'h00000000 /* 0x27cc */;
                2548: data_o = 32'h00000000 /* 0x27d0 */;
                2549: data_o = 32'h00000000 /* 0x27d4 */;
                2550: data_o = 32'h00000000 /* 0x27d8 */;
                2551: data_o = 32'h00000000 /* 0x27dc */;
                2552: data_o = 32'h00000000 /* 0x27e0 */;
                2553: data_o = 32'h00000000 /* 0x27e4 */;
                2554: data_o = 32'h00000000 /* 0x27e8 */;
                2555: data_o = 32'h00000000 /* 0x27ec */;
                2556: data_o = 32'h00000000 /* 0x27f0 */;
                2557: data_o = 32'h00000000 /* 0x27f4 */;
                2558: data_o = 32'h00000000 /* 0x27f8 */;
                2559: data_o = 32'h00000000 /* 0x27fc */;
                2560: data_o = 32'h00000000 /* 0x2800 */;
                2561: data_o = 32'h00000000 /* 0x2804 */;
                2562: data_o = 32'h00000000 /* 0x2808 */;
                2563: data_o = 32'h00000000 /* 0x280c */;
                2564: data_o = 32'h00000000 /* 0x2810 */;
                2565: data_o = 32'h00000000 /* 0x2814 */;
                2566: data_o = 32'h00000000 /* 0x2818 */;
                2567: data_o = 32'h00000000 /* 0x281c */;
                2568: data_o = 32'h00000000 /* 0x2820 */;
                2569: data_o = 32'h00000000 /* 0x2824 */;
                2570: data_o = 32'h00000000 /* 0x2828 */;
                2571: data_o = 32'h00000000 /* 0x282c */;
                2572: data_o = 32'h00000000 /* 0x2830 */;
                2573: data_o = 32'h00000000 /* 0x2834 */;
                2574: data_o = 32'h00000000 /* 0x2838 */;
                2575: data_o = 32'h00000000 /* 0x283c */;
                2576: data_o = 32'h00000000 /* 0x2840 */;
                2577: data_o = 32'h00000000 /* 0x2844 */;
                2578: data_o = 32'h00000000 /* 0x2848 */;
                2579: data_o = 32'h00000000 /* 0x284c */;
                2580: data_o = 32'h00000000 /* 0x2850 */;
                2581: data_o = 32'h00000000 /* 0x2854 */;
                2582: data_o = 32'h00000000 /* 0x2858 */;
                2583: data_o = 32'h00000000 /* 0x285c */;
                2584: data_o = 32'h00000000 /* 0x2860 */;
                2585: data_o = 32'h00000000 /* 0x2864 */;
                2586: data_o = 32'h00000000 /* 0x2868 */;
                2587: data_o = 32'h00000000 /* 0x286c */;
                2588: data_o = 32'h00000000 /* 0x2870 */;
                2589: data_o = 32'h00000000 /* 0x2874 */;
                2590: data_o = 32'h00000000 /* 0x2878 */;
                2591: data_o = 32'h00000000 /* 0x287c */;
                2592: data_o = 32'h00000000 /* 0x2880 */;
                2593: data_o = 32'h00000000 /* 0x2884 */;
                2594: data_o = 32'h00000000 /* 0x2888 */;
                2595: data_o = 32'h00000000 /* 0x288c */;
                2596: data_o = 32'h00000000 /* 0x2890 */;
                2597: data_o = 32'h00000000 /* 0x2894 */;
                2598: data_o = 32'h00000000 /* 0x2898 */;
                2599: data_o = 32'h00000000 /* 0x289c */;
                2600: data_o = 32'h00000000 /* 0x28a0 */;
                2601: data_o = 32'h00000000 /* 0x28a4 */;
                2602: data_o = 32'h00000000 /* 0x28a8 */;
                2603: data_o = 32'h00000000 /* 0x28ac */;
                2604: data_o = 32'h00000000 /* 0x28b0 */;
                2605: data_o = 32'h00000000 /* 0x28b4 */;
                2606: data_o = 32'h00000000 /* 0x28b8 */;
                2607: data_o = 32'h00000000 /* 0x28bc */;
                2608: data_o = 32'h00000000 /* 0x28c0 */;
                2609: data_o = 32'h00000000 /* 0x28c4 */;
                2610: data_o = 32'h00000000 /* 0x28c8 */;
                2611: data_o = 32'h00000000 /* 0x28cc */;
                2612: data_o = 32'h00000000 /* 0x28d0 */;
                2613: data_o = 32'h00000000 /* 0x28d4 */;
                2614: data_o = 32'h00000000 /* 0x28d8 */;
                2615: data_o = 32'h00000000 /* 0x28dc */;
                2616: data_o = 32'h00000000 /* 0x28e0 */;
                2617: data_o = 32'h00000000 /* 0x28e4 */;
                2618: data_o = 32'h00000000 /* 0x28e8 */;
                2619: data_o = 32'h00000000 /* 0x28ec */;
                2620: data_o = 32'h00000000 /* 0x28f0 */;
                2621: data_o = 32'h00000000 /* 0x28f4 */;
                2622: data_o = 32'h00000000 /* 0x28f8 */;
                2623: data_o = 32'h00000000 /* 0x28fc */;
                2624: data_o = 32'h00000000 /* 0x2900 */;
                2625: data_o = 32'h00000000 /* 0x2904 */;
                2626: data_o = 32'h00000000 /* 0x2908 */;
                2627: data_o = 32'h00000000 /* 0x290c */;
                2628: data_o = 32'h00000000 /* 0x2910 */;
                2629: data_o = 32'h00000000 /* 0x2914 */;
                2630: data_o = 32'h00000000 /* 0x2918 */;
                2631: data_o = 32'h00000000 /* 0x291c */;
                2632: data_o = 32'h00000000 /* 0x2920 */;
                2633: data_o = 32'h00000000 /* 0x2924 */;
                2634: data_o = 32'h00000000 /* 0x2928 */;
                2635: data_o = 32'h00000000 /* 0x292c */;
                2636: data_o = 32'h00000000 /* 0x2930 */;
                2637: data_o = 32'h00000000 /* 0x2934 */;
                2638: data_o = 32'h00000000 /* 0x2938 */;
                2639: data_o = 32'h00000000 /* 0x293c */;
                2640: data_o = 32'h00000000 /* 0x2940 */;
                2641: data_o = 32'h00000000 /* 0x2944 */;
                2642: data_o = 32'h00000000 /* 0x2948 */;
                2643: data_o = 32'h00000000 /* 0x294c */;
                2644: data_o = 32'h00000000 /* 0x2950 */;
                2645: data_o = 32'h00000000 /* 0x2954 */;
                2646: data_o = 32'h00000000 /* 0x2958 */;
                2647: data_o = 32'h00000000 /* 0x295c */;
                2648: data_o = 32'h00000000 /* 0x2960 */;
                2649: data_o = 32'h00000000 /* 0x2964 */;
                2650: data_o = 32'h00000000 /* 0x2968 */;
                2651: data_o = 32'h00000000 /* 0x296c */;
                2652: data_o = 32'h00000000 /* 0x2970 */;
                2653: data_o = 32'h00000000 /* 0x2974 */;
                2654: data_o = 32'h00000000 /* 0x2978 */;
                2655: data_o = 32'h00000000 /* 0x297c */;
                2656: data_o = 32'h00000000 /* 0x2980 */;
                2657: data_o = 32'h00000000 /* 0x2984 */;
                2658: data_o = 32'h00000000 /* 0x2988 */;
                2659: data_o = 32'h00000000 /* 0x298c */;
                2660: data_o = 32'h00000000 /* 0x2990 */;
                2661: data_o = 32'h00000000 /* 0x2994 */;
                2662: data_o = 32'h00000000 /* 0x2998 */;
                2663: data_o = 32'h00000000 /* 0x299c */;
                2664: data_o = 32'h00000000 /* 0x29a0 */;
                2665: data_o = 32'h00000000 /* 0x29a4 */;
                2666: data_o = 32'h00000000 /* 0x29a8 */;
                2667: data_o = 32'h00000000 /* 0x29ac */;
                2668: data_o = 32'h00000000 /* 0x29b0 */;
                2669: data_o = 32'h00000000 /* 0x29b4 */;
                2670: data_o = 32'h00000000 /* 0x29b8 */;
                2671: data_o = 32'h00000000 /* 0x29bc */;
                2672: data_o = 32'h00000000 /* 0x29c0 */;
                2673: data_o = 32'h00000000 /* 0x29c4 */;
                2674: data_o = 32'h00000000 /* 0x29c8 */;
                2675: data_o = 32'h00000000 /* 0x29cc */;
                2676: data_o = 32'h00000000 /* 0x29d0 */;
                2677: data_o = 32'h00000000 /* 0x29d4 */;
                2678: data_o = 32'h00000000 /* 0x29d8 */;
                2679: data_o = 32'h00000000 /* 0x29dc */;
                2680: data_o = 32'h00000000 /* 0x29e0 */;
                2681: data_o = 32'h00000000 /* 0x29e4 */;
                2682: data_o = 32'h00000000 /* 0x29e8 */;
                2683: data_o = 32'h00000000 /* 0x29ec */;
                2684: data_o = 32'h00000000 /* 0x29f0 */;
                2685: data_o = 32'h00000000 /* 0x29f4 */;
                2686: data_o = 32'h00000000 /* 0x29f8 */;
                2687: data_o = 32'h00000000 /* 0x29fc */;
                2688: data_o = 32'h00000000 /* 0x2a00 */;
                2689: data_o = 32'h00000000 /* 0x2a04 */;
                2690: data_o = 32'h00000000 /* 0x2a08 */;
                2691: data_o = 32'h00000000 /* 0x2a0c */;
                2692: data_o = 32'h00000000 /* 0x2a10 */;
                2693: data_o = 32'h00000000 /* 0x2a14 */;
                2694: data_o = 32'h00000000 /* 0x2a18 */;
                2695: data_o = 32'h00000000 /* 0x2a1c */;
                2696: data_o = 32'h00000000 /* 0x2a20 */;
                2697: data_o = 32'h00000000 /* 0x2a24 */;
                2698: data_o = 32'h00000000 /* 0x2a28 */;
                2699: data_o = 32'h00000000 /* 0x2a2c */;
                2700: data_o = 32'h00000000 /* 0x2a30 */;
                2701: data_o = 32'h00000000 /* 0x2a34 */;
                2702: data_o = 32'h00000000 /* 0x2a38 */;
                2703: data_o = 32'h00000000 /* 0x2a3c */;
                2704: data_o = 32'h00000000 /* 0x2a40 */;
                2705: data_o = 32'h00000000 /* 0x2a44 */;
                2706: data_o = 32'h00000000 /* 0x2a48 */;
                2707: data_o = 32'h00000000 /* 0x2a4c */;
                2708: data_o = 32'h00000000 /* 0x2a50 */;
                2709: data_o = 32'h00000000 /* 0x2a54 */;
                2710: data_o = 32'h00000000 /* 0x2a58 */;
                2711: data_o = 32'h00000000 /* 0x2a5c */;
                2712: data_o = 32'h00000000 /* 0x2a60 */;
                2713: data_o = 32'h00000000 /* 0x2a64 */;
                2714: data_o = 32'h00000000 /* 0x2a68 */;
                2715: data_o = 32'h00000000 /* 0x2a6c */;
                2716: data_o = 32'h00000000 /* 0x2a70 */;
                2717: data_o = 32'h00000000 /* 0x2a74 */;
                2718: data_o = 32'h00000000 /* 0x2a78 */;
                2719: data_o = 32'h00000000 /* 0x2a7c */;
                2720: data_o = 32'h00000000 /* 0x2a80 */;
                2721: data_o = 32'h00000000 /* 0x2a84 */;
                2722: data_o = 32'h00000000 /* 0x2a88 */;
                2723: data_o = 32'h00000000 /* 0x2a8c */;
                2724: data_o = 32'h00000000 /* 0x2a90 */;
                2725: data_o = 32'h00000000 /* 0x2a94 */;
                2726: data_o = 32'h00000000 /* 0x2a98 */;
                2727: data_o = 32'h00000000 /* 0x2a9c */;
                2728: data_o = 32'h00000000 /* 0x2aa0 */;
                2729: data_o = 32'h00000000 /* 0x2aa4 */;
                2730: data_o = 32'h00000000 /* 0x2aa8 */;
                2731: data_o = 32'h00000000 /* 0x2aac */;
                2732: data_o = 32'h00000000 /* 0x2ab0 */;
                2733: data_o = 32'h00000000 /* 0x2ab4 */;
                2734: data_o = 32'h00000000 /* 0x2ab8 */;
                2735: data_o = 32'h00000000 /* 0x2abc */;
                2736: data_o = 32'h00000000 /* 0x2ac0 */;
                2737: data_o = 32'h00000000 /* 0x2ac4 */;
                2738: data_o = 32'h00000000 /* 0x2ac8 */;
                2739: data_o = 32'h00000000 /* 0x2acc */;
                2740: data_o = 32'h00000000 /* 0x2ad0 */;
                2741: data_o = 32'h00000000 /* 0x2ad4 */;
                2742: data_o = 32'h00000000 /* 0x2ad8 */;
                2743: data_o = 32'h00000000 /* 0x2adc */;
                2744: data_o = 32'h00000000 /* 0x2ae0 */;
                2745: data_o = 32'h00000000 /* 0x2ae4 */;
                2746: data_o = 32'h00000000 /* 0x2ae8 */;
                2747: data_o = 32'h00000000 /* 0x2aec */;
                2748: data_o = 32'h00000000 /* 0x2af0 */;
                2749: data_o = 32'h00000000 /* 0x2af4 */;
                2750: data_o = 32'h00000000 /* 0x2af8 */;
                2751: data_o = 32'h00000000 /* 0x2afc */;
                2752: data_o = 32'h00000000 /* 0x2b00 */;
                2753: data_o = 32'h00000000 /* 0x2b04 */;
                2754: data_o = 32'h00000000 /* 0x2b08 */;
                2755: data_o = 32'h00000000 /* 0x2b0c */;
                2756: data_o = 32'h00000000 /* 0x2b10 */;
                2757: data_o = 32'h00000000 /* 0x2b14 */;
                2758: data_o = 32'h00000000 /* 0x2b18 */;
                2759: data_o = 32'h00000000 /* 0x2b1c */;
                2760: data_o = 32'h00000000 /* 0x2b20 */;
                2761: data_o = 32'h00000000 /* 0x2b24 */;
                2762: data_o = 32'h00000000 /* 0x2b28 */;
                2763: data_o = 32'h00000000 /* 0x2b2c */;
                2764: data_o = 32'h00000000 /* 0x2b30 */;
                2765: data_o = 32'h00000000 /* 0x2b34 */;
                2766: data_o = 32'h00000000 /* 0x2b38 */;
                2767: data_o = 32'h00000000 /* 0x2b3c */;
                2768: data_o = 32'h00000000 /* 0x2b40 */;
                2769: data_o = 32'h00000000 /* 0x2b44 */;
                2770: data_o = 32'h00000000 /* 0x2b48 */;
                2771: data_o = 32'h00000000 /* 0x2b4c */;
                2772: data_o = 32'h00000000 /* 0x2b50 */;
                2773: data_o = 32'h00000000 /* 0x2b54 */;
                2774: data_o = 32'h00000000 /* 0x2b58 */;
                2775: data_o = 32'h00000000 /* 0x2b5c */;
                2776: data_o = 32'h00000000 /* 0x2b60 */;
                2777: data_o = 32'h00000000 /* 0x2b64 */;
                2778: data_o = 32'h00000000 /* 0x2b68 */;
                2779: data_o = 32'h00000000 /* 0x2b6c */;
                2780: data_o = 32'h00000000 /* 0x2b70 */;
                2781: data_o = 32'h00000000 /* 0x2b74 */;
                2782: data_o = 32'h00000000 /* 0x2b78 */;
                2783: data_o = 32'h00000000 /* 0x2b7c */;
                2784: data_o = 32'h00000000 /* 0x2b80 */;
                2785: data_o = 32'h00000000 /* 0x2b84 */;
                2786: data_o = 32'h00000000 /* 0x2b88 */;
                2787: data_o = 32'h00000000 /* 0x2b8c */;
                2788: data_o = 32'h00000000 /* 0x2b90 */;
                2789: data_o = 32'h00000000 /* 0x2b94 */;
                2790: data_o = 32'h00000000 /* 0x2b98 */;
                2791: data_o = 32'h00000000 /* 0x2b9c */;
                2792: data_o = 32'h00000000 /* 0x2ba0 */;
                2793: data_o = 32'h00000000 /* 0x2ba4 */;
                2794: data_o = 32'h00000000 /* 0x2ba8 */;
                2795: data_o = 32'h00000000 /* 0x2bac */;
                2796: data_o = 32'h00000000 /* 0x2bb0 */;
                2797: data_o = 32'h00000000 /* 0x2bb4 */;
                2798: data_o = 32'h00000000 /* 0x2bb8 */;
                2799: data_o = 32'h00000000 /* 0x2bbc */;
                2800: data_o = 32'h00000000 /* 0x2bc0 */;
                2801: data_o = 32'h00000000 /* 0x2bc4 */;
                2802: data_o = 32'h00000000 /* 0x2bc8 */;
                2803: data_o = 32'h00000000 /* 0x2bcc */;
                2804: data_o = 32'h00000000 /* 0x2bd0 */;
                2805: data_o = 32'h00000000 /* 0x2bd4 */;
                2806: data_o = 32'h00000000 /* 0x2bd8 */;
                2807: data_o = 32'h00000000 /* 0x2bdc */;
                2808: data_o = 32'h00000000 /* 0x2be0 */;
                2809: data_o = 32'h00000000 /* 0x2be4 */;
                2810: data_o = 32'h00000000 /* 0x2be8 */;
                2811: data_o = 32'h00000000 /* 0x2bec */;
                2812: data_o = 32'h00000000 /* 0x2bf0 */;
                2813: data_o = 32'h00000000 /* 0x2bf4 */;
                2814: data_o = 32'h00000000 /* 0x2bf8 */;
                2815: data_o = 32'h00000000 /* 0x2bfc */;
                2816: data_o = 32'h00000000 /* 0x2c00 */;
                2817: data_o = 32'h00000000 /* 0x2c04 */;
                2818: data_o = 32'h00000000 /* 0x2c08 */;
                2819: data_o = 32'h00000000 /* 0x2c0c */;
                2820: data_o = 32'h00000000 /* 0x2c10 */;
                2821: data_o = 32'h00000000 /* 0x2c14 */;
                2822: data_o = 32'h00000000 /* 0x2c18 */;
                2823: data_o = 32'h00000000 /* 0x2c1c */;
                2824: data_o = 32'h00000000 /* 0x2c20 */;
                2825: data_o = 32'h00000000 /* 0x2c24 */;
                2826: data_o = 32'h00000000 /* 0x2c28 */;
                2827: data_o = 32'h00000000 /* 0x2c2c */;
                2828: data_o = 32'h00000000 /* 0x2c30 */;
                2829: data_o = 32'h00000000 /* 0x2c34 */;
                2830: data_o = 32'h00000000 /* 0x2c38 */;
                2831: data_o = 32'h00000000 /* 0x2c3c */;
                2832: data_o = 32'h00000000 /* 0x2c40 */;
                2833: data_o = 32'h00000000 /* 0x2c44 */;
                2834: data_o = 32'h00000000 /* 0x2c48 */;
                2835: data_o = 32'h00000000 /* 0x2c4c */;
                2836: data_o = 32'h00000000 /* 0x2c50 */;
                2837: data_o = 32'h00000000 /* 0x2c54 */;
                2838: data_o = 32'h00000000 /* 0x2c58 */;
                2839: data_o = 32'h00000000 /* 0x2c5c */;
                2840: data_o = 32'h00000000 /* 0x2c60 */;
                2841: data_o = 32'h00000000 /* 0x2c64 */;
                2842: data_o = 32'h00000000 /* 0x2c68 */;
                2843: data_o = 32'h00000000 /* 0x2c6c */;
                2844: data_o = 32'h00000000 /* 0x2c70 */;
                2845: data_o = 32'h00000000 /* 0x2c74 */;
                2846: data_o = 32'h00000000 /* 0x2c78 */;
                2847: data_o = 32'h00000000 /* 0x2c7c */;
                2848: data_o = 32'h00000000 /* 0x2c80 */;
                2849: data_o = 32'h00000000 /* 0x2c84 */;
                2850: data_o = 32'h00000000 /* 0x2c88 */;
                2851: data_o = 32'h00000000 /* 0x2c8c */;
                2852: data_o = 32'h00000000 /* 0x2c90 */;
                2853: data_o = 32'h00000000 /* 0x2c94 */;
                2854: data_o = 32'h00000000 /* 0x2c98 */;
                2855: data_o = 32'h00000000 /* 0x2c9c */;
                2856: data_o = 32'h00000000 /* 0x2ca0 */;
                2857: data_o = 32'h00000000 /* 0x2ca4 */;
                2858: data_o = 32'h00000000 /* 0x2ca8 */;
                2859: data_o = 32'h00000000 /* 0x2cac */;
                2860: data_o = 32'h00000000 /* 0x2cb0 */;
                2861: data_o = 32'h00000000 /* 0x2cb4 */;
                2862: data_o = 32'h00000000 /* 0x2cb8 */;
                2863: data_o = 32'h00000000 /* 0x2cbc */;
                2864: data_o = 32'h00000000 /* 0x2cc0 */;
                2865: data_o = 32'h00000000 /* 0x2cc4 */;
                2866: data_o = 32'h00000000 /* 0x2cc8 */;
                2867: data_o = 32'h00000000 /* 0x2ccc */;
                2868: data_o = 32'h00000000 /* 0x2cd0 */;
                2869: data_o = 32'h00000000 /* 0x2cd4 */;
                2870: data_o = 32'h00000000 /* 0x2cd8 */;
                2871: data_o = 32'h00000000 /* 0x2cdc */;
                2872: data_o = 32'h00000000 /* 0x2ce0 */;
                2873: data_o = 32'h00000000 /* 0x2ce4 */;
                2874: data_o = 32'h00000000 /* 0x2ce8 */;
                2875: data_o = 32'h00000000 /* 0x2cec */;
                2876: data_o = 32'h00000000 /* 0x2cf0 */;
                2877: data_o = 32'h00000000 /* 0x2cf4 */;
                2878: data_o = 32'h00000000 /* 0x2cf8 */;
                2879: data_o = 32'h00000000 /* 0x2cfc */;
                2880: data_o = 32'h00000000 /* 0x2d00 */;
                2881: data_o = 32'h00000000 /* 0x2d04 */;
                2882: data_o = 32'h00000000 /* 0x2d08 */;
                2883: data_o = 32'h00000000 /* 0x2d0c */;
                2884: data_o = 32'h00000000 /* 0x2d10 */;
                2885: data_o = 32'h00000000 /* 0x2d14 */;
                2886: data_o = 32'h00000000 /* 0x2d18 */;
                2887: data_o = 32'h00000000 /* 0x2d1c */;
                2888: data_o = 32'h00000000 /* 0x2d20 */;
                2889: data_o = 32'h00000000 /* 0x2d24 */;
                2890: data_o = 32'h00000000 /* 0x2d28 */;
                2891: data_o = 32'h00000000 /* 0x2d2c */;
                2892: data_o = 32'h00000000 /* 0x2d30 */;
                2893: data_o = 32'h00000000 /* 0x2d34 */;
                2894: data_o = 32'h00000000 /* 0x2d38 */;
                2895: data_o = 32'h00000000 /* 0x2d3c */;
                2896: data_o = 32'h00000000 /* 0x2d40 */;
                2897: data_o = 32'h00000000 /* 0x2d44 */;
                2898: data_o = 32'h00000000 /* 0x2d48 */;
                2899: data_o = 32'h00000000 /* 0x2d4c */;
                2900: data_o = 32'h00000000 /* 0x2d50 */;
                2901: data_o = 32'h00000000 /* 0x2d54 */;
                2902: data_o = 32'h00000000 /* 0x2d58 */;
                2903: data_o = 32'h00000000 /* 0x2d5c */;
                2904: data_o = 32'h00000000 /* 0x2d60 */;
                2905: data_o = 32'h00000000 /* 0x2d64 */;
                2906: data_o = 32'h00000000 /* 0x2d68 */;
                2907: data_o = 32'h00000000 /* 0x2d6c */;
                2908: data_o = 32'h00000000 /* 0x2d70 */;
                2909: data_o = 32'h00000000 /* 0x2d74 */;
                2910: data_o = 32'h00000000 /* 0x2d78 */;
                2911: data_o = 32'h00000000 /* 0x2d7c */;
                2912: data_o = 32'h00000000 /* 0x2d80 */;
                2913: data_o = 32'h00000000 /* 0x2d84 */;
                2914: data_o = 32'h00000000 /* 0x2d88 */;
                2915: data_o = 32'h00000000 /* 0x2d8c */;
                2916: data_o = 32'h00000000 /* 0x2d90 */;
                2917: data_o = 32'h00000000 /* 0x2d94 */;
                2918: data_o = 32'h00000000 /* 0x2d98 */;
                2919: data_o = 32'h00000000 /* 0x2d9c */;
                2920: data_o = 32'h00000000 /* 0x2da0 */;
                2921: data_o = 32'h00000000 /* 0x2da4 */;
                2922: data_o = 32'h00000000 /* 0x2da8 */;
                2923: data_o = 32'h00000000 /* 0x2dac */;
                2924: data_o = 32'h00000000 /* 0x2db0 */;
                2925: data_o = 32'h00000000 /* 0x2db4 */;
                2926: data_o = 32'h00000000 /* 0x2db8 */;
                2927: data_o = 32'h00000000 /* 0x2dbc */;
                2928: data_o = 32'h00000000 /* 0x2dc0 */;
                2929: data_o = 32'h00000000 /* 0x2dc4 */;
                2930: data_o = 32'h00000000 /* 0x2dc8 */;
                2931: data_o = 32'h00000000 /* 0x2dcc */;
                2932: data_o = 32'h00000000 /* 0x2dd0 */;
                2933: data_o = 32'h00000000 /* 0x2dd4 */;
                2934: data_o = 32'h00000000 /* 0x2dd8 */;
                2935: data_o = 32'h00000000 /* 0x2ddc */;
                2936: data_o = 32'h00000000 /* 0x2de0 */;
                2937: data_o = 32'h00000000 /* 0x2de4 */;
                2938: data_o = 32'h00000000 /* 0x2de8 */;
                2939: data_o = 32'h00000000 /* 0x2dec */;
                2940: data_o = 32'h00000000 /* 0x2df0 */;
                2941: data_o = 32'h00000000 /* 0x2df4 */;
                2942: data_o = 32'h00000000 /* 0x2df8 */;
                2943: data_o = 32'h00000000 /* 0x2dfc */;
                2944: data_o = 32'h00000000 /* 0x2e00 */;
                2945: data_o = 32'h00000000 /* 0x2e04 */;
                2946: data_o = 32'h00000000 /* 0x2e08 */;
                2947: data_o = 32'h00000000 /* 0x2e0c */;
                2948: data_o = 32'h00000000 /* 0x2e10 */;
                2949: data_o = 32'h00000000 /* 0x2e14 */;
                2950: data_o = 32'h00000000 /* 0x2e18 */;
                2951: data_o = 32'h00000000 /* 0x2e1c */;
                2952: data_o = 32'h00000000 /* 0x2e20 */;
                2953: data_o = 32'h00000000 /* 0x2e24 */;
                2954: data_o = 32'h00000000 /* 0x2e28 */;
                2955: data_o = 32'h00000000 /* 0x2e2c */;
                2956: data_o = 32'h00000000 /* 0x2e30 */;
                2957: data_o = 32'h00000000 /* 0x2e34 */;
                2958: data_o = 32'h00000000 /* 0x2e38 */;
                2959: data_o = 32'h00000000 /* 0x2e3c */;
                2960: data_o = 32'h00000000 /* 0x2e40 */;
                2961: data_o = 32'h00000000 /* 0x2e44 */;
                2962: data_o = 32'h00000000 /* 0x2e48 */;
                2963: data_o = 32'h00000000 /* 0x2e4c */;
                2964: data_o = 32'h00000000 /* 0x2e50 */;
                2965: data_o = 32'h00000000 /* 0x2e54 */;
                2966: data_o = 32'h00000000 /* 0x2e58 */;
                2967: data_o = 32'h00000000 /* 0x2e5c */;
                2968: data_o = 32'h00000000 /* 0x2e60 */;
                2969: data_o = 32'h00000000 /* 0x2e64 */;
                2970: data_o = 32'h00000000 /* 0x2e68 */;
                2971: data_o = 32'h00000000 /* 0x2e6c */;
                2972: data_o = 32'h00000000 /* 0x2e70 */;
                2973: data_o = 32'h00000000 /* 0x2e74 */;
                2974: data_o = 32'h00000000 /* 0x2e78 */;
                2975: data_o = 32'h00000000 /* 0x2e7c */;
                2976: data_o = 32'h00000000 /* 0x2e80 */;
                2977: data_o = 32'h00000000 /* 0x2e84 */;
                2978: data_o = 32'h00000000 /* 0x2e88 */;
                2979: data_o = 32'h00000000 /* 0x2e8c */;
                2980: data_o = 32'h00000000 /* 0x2e90 */;
                2981: data_o = 32'h00000000 /* 0x2e94 */;
                2982: data_o = 32'h00000000 /* 0x2e98 */;
                2983: data_o = 32'h00000000 /* 0x2e9c */;
                2984: data_o = 32'h00000000 /* 0x2ea0 */;
                2985: data_o = 32'h00000000 /* 0x2ea4 */;
                2986: data_o = 32'h00000000 /* 0x2ea8 */;
                2987: data_o = 32'h00000000 /* 0x2eac */;
                2988: data_o = 32'h00000000 /* 0x2eb0 */;
                2989: data_o = 32'h00000000 /* 0x2eb4 */;
                2990: data_o = 32'h00000000 /* 0x2eb8 */;
                2991: data_o = 32'h00000000 /* 0x2ebc */;
                2992: data_o = 32'h00000000 /* 0x2ec0 */;
                2993: data_o = 32'h00000000 /* 0x2ec4 */;
                2994: data_o = 32'h00000000 /* 0x2ec8 */;
                2995: data_o = 32'h00000000 /* 0x2ecc */;
                2996: data_o = 32'h00000000 /* 0x2ed0 */;
                2997: data_o = 32'h00000000 /* 0x2ed4 */;
                2998: data_o = 32'h00000000 /* 0x2ed8 */;
                2999: data_o = 32'h00000000 /* 0x2edc */;
                3000: data_o = 32'h00000000 /* 0x2ee0 */;
                3001: data_o = 32'h00000000 /* 0x2ee4 */;
                3002: data_o = 32'h00000000 /* 0x2ee8 */;
                3003: data_o = 32'h00000000 /* 0x2eec */;
                3004: data_o = 32'h00000000 /* 0x2ef0 */;
                3005: data_o = 32'h00000000 /* 0x2ef4 */;
                3006: data_o = 32'h00000000 /* 0x2ef8 */;
                3007: data_o = 32'h00000000 /* 0x2efc */;
                3008: data_o = 32'h00000000 /* 0x2f00 */;
                3009: data_o = 32'h00000000 /* 0x2f04 */;
                3010: data_o = 32'h00000000 /* 0x2f08 */;
                3011: data_o = 32'h00000000 /* 0x2f0c */;
                3012: data_o = 32'h00000000 /* 0x2f10 */;
                3013: data_o = 32'h00000000 /* 0x2f14 */;
                3014: data_o = 32'h00000000 /* 0x2f18 */;
                3015: data_o = 32'h00000000 /* 0x2f1c */;
                3016: data_o = 32'h00000000 /* 0x2f20 */;
                3017: data_o = 32'h00000000 /* 0x2f24 */;
                3018: data_o = 32'h00000000 /* 0x2f28 */;
                3019: data_o = 32'h00000000 /* 0x2f2c */;
                3020: data_o = 32'h00000000 /* 0x2f30 */;
                3021: data_o = 32'h00000000 /* 0x2f34 */;
                3022: data_o = 32'h00000000 /* 0x2f38 */;
                3023: data_o = 32'h00000000 /* 0x2f3c */;
                3024: data_o = 32'h00000000 /* 0x2f40 */;
                3025: data_o = 32'h00000000 /* 0x2f44 */;
                3026: data_o = 32'h00000000 /* 0x2f48 */;
                3027: data_o = 32'h00000000 /* 0x2f4c */;
                3028: data_o = 32'h00000000 /* 0x2f50 */;
                3029: data_o = 32'h00000000 /* 0x2f54 */;
                3030: data_o = 32'h00000000 /* 0x2f58 */;
                3031: data_o = 32'h00000000 /* 0x2f5c */;
                3032: data_o = 32'h00000000 /* 0x2f60 */;
                3033: data_o = 32'h00000000 /* 0x2f64 */;
                3034: data_o = 32'h00000000 /* 0x2f68 */;
                3035: data_o = 32'h00000000 /* 0x2f6c */;
                3036: data_o = 32'h00000000 /* 0x2f70 */;
                3037: data_o = 32'h00000000 /* 0x2f74 */;
                3038: data_o = 32'h00000000 /* 0x2f78 */;
                3039: data_o = 32'h00000000 /* 0x2f7c */;
                3040: data_o = 32'h00000000 /* 0x2f80 */;
                3041: data_o = 32'h00000000 /* 0x2f84 */;
                3042: data_o = 32'h00000000 /* 0x2f88 */;
                3043: data_o = 32'h00000000 /* 0x2f8c */;
                3044: data_o = 32'h00000000 /* 0x2f90 */;
                3045: data_o = 32'h00000000 /* 0x2f94 */;
                3046: data_o = 32'h00000000 /* 0x2f98 */;
                3047: data_o = 32'h00000000 /* 0x2f9c */;
                3048: data_o = 32'h00000000 /* 0x2fa0 */;
                3049: data_o = 32'h00000000 /* 0x2fa4 */;
                3050: data_o = 32'h00000000 /* 0x2fa8 */;
                3051: data_o = 32'h00000000 /* 0x2fac */;
                3052: data_o = 32'h00000000 /* 0x2fb0 */;
                3053: data_o = 32'h00000000 /* 0x2fb4 */;
                3054: data_o = 32'h00000000 /* 0x2fb8 */;
                3055: data_o = 32'h00000000 /* 0x2fbc */;
                3056: data_o = 32'h00000000 /* 0x2fc0 */;
                3057: data_o = 32'h00000000 /* 0x2fc4 */;
                3058: data_o = 32'h00000000 /* 0x2fc8 */;
                3059: data_o = 32'h00000000 /* 0x2fcc */;
                3060: data_o = 32'h00000000 /* 0x2fd0 */;
                3061: data_o = 32'h00000000 /* 0x2fd4 */;
                3062: data_o = 32'h00000000 /* 0x2fd8 */;
                3063: data_o = 32'h00000000 /* 0x2fdc */;
                3064: data_o = 32'h00000000 /* 0x2fe0 */;
                3065: data_o = 32'h00000000 /* 0x2fe4 */;
                3066: data_o = 32'h00000000 /* 0x2fe8 */;
                3067: data_o = 32'h00000000 /* 0x2fec */;
                3068: data_o = 32'h00000000 /* 0x2ff0 */;
                3069: data_o = 32'h00000000 /* 0x2ff4 */;
                3070: data_o = 32'h00000000 /* 0x2ff8 */;
                3071: data_o = 32'h00000000 /* 0x2ffc */;
                3072: data_o = 32'h00000000 /* 0x3000 */;
                3073: data_o = 32'h00000000 /* 0x3004 */;
                3074: data_o = 32'h00000000 /* 0x3008 */;
                3075: data_o = 32'h00000000 /* 0x300c */;
                3076: data_o = 32'h00000000 /* 0x3010 */;
                3077: data_o = 32'h00000000 /* 0x3014 */;
                3078: data_o = 32'h00000000 /* 0x3018 */;
                3079: data_o = 32'h00000000 /* 0x301c */;
                3080: data_o = 32'h00000000 /* 0x3020 */;
                3081: data_o = 32'h00000000 /* 0x3024 */;
                3082: data_o = 32'h00000000 /* 0x3028 */;
                3083: data_o = 32'h00000000 /* 0x302c */;
                3084: data_o = 32'h00000000 /* 0x3030 */;
                3085: data_o = 32'h00000000 /* 0x3034 */;
                3086: data_o = 32'h00000000 /* 0x3038 */;
                3087: data_o = 32'h00000000 /* 0x303c */;
                3088: data_o = 32'h00000000 /* 0x3040 */;
                3089: data_o = 32'h00000000 /* 0x3044 */;
                3090: data_o = 32'h00000000 /* 0x3048 */;
                3091: data_o = 32'h00000000 /* 0x304c */;
                3092: data_o = 32'h00000000 /* 0x3050 */;
                3093: data_o = 32'h00000000 /* 0x3054 */;
                3094: data_o = 32'h00000000 /* 0x3058 */;
                3095: data_o = 32'h00000000 /* 0x305c */;
                3096: data_o = 32'h00000000 /* 0x3060 */;
                3097: data_o = 32'h00000000 /* 0x3064 */;
                3098: data_o = 32'h00000000 /* 0x3068 */;
                3099: data_o = 32'h00000000 /* 0x306c */;
                3100: data_o = 32'h00000000 /* 0x3070 */;
                3101: data_o = 32'h00000000 /* 0x3074 */;
                3102: data_o = 32'h00000000 /* 0x3078 */;
                3103: data_o = 32'h00000000 /* 0x307c */;
                3104: data_o = 32'h00000000 /* 0x3080 */;
                3105: data_o = 32'h00000000 /* 0x3084 */;
                3106: data_o = 32'h00000000 /* 0x3088 */;
                3107: data_o = 32'h00000000 /* 0x308c */;
                3108: data_o = 32'h00000000 /* 0x3090 */;
                3109: data_o = 32'h00000000 /* 0x3094 */;
                3110: data_o = 32'h00000000 /* 0x3098 */;
                3111: data_o = 32'h00000000 /* 0x309c */;
                3112: data_o = 32'h00000000 /* 0x30a0 */;
                3113: data_o = 32'h00000000 /* 0x30a4 */;
                3114: data_o = 32'h00000000 /* 0x30a8 */;
                3115: data_o = 32'h00000000 /* 0x30ac */;
                3116: data_o = 32'h00000000 /* 0x30b0 */;
                3117: data_o = 32'h00000000 /* 0x30b4 */;
                3118: data_o = 32'h00000000 /* 0x30b8 */;
                3119: data_o = 32'h00000000 /* 0x30bc */;
                3120: data_o = 32'h00000000 /* 0x30c0 */;
                3121: data_o = 32'h00000000 /* 0x30c4 */;
                3122: data_o = 32'h00000000 /* 0x30c8 */;
                3123: data_o = 32'h00000000 /* 0x30cc */;
                3124: data_o = 32'h00000000 /* 0x30d0 */;
                3125: data_o = 32'h00000000 /* 0x30d4 */;
                3126: data_o = 32'h00000000 /* 0x30d8 */;
                3127: data_o = 32'h00000000 /* 0x30dc */;
                3128: data_o = 32'h00000000 /* 0x30e0 */;
                3129: data_o = 32'h00000000 /* 0x30e4 */;
                3130: data_o = 32'h00000000 /* 0x30e8 */;
                3131: data_o = 32'h00000000 /* 0x30ec */;
                3132: data_o = 32'h00000000 /* 0x30f0 */;
                3133: data_o = 32'h00000000 /* 0x30f4 */;
                3134: data_o = 32'h00000000 /* 0x30f8 */;
                3135: data_o = 32'h00000000 /* 0x30fc */;
                3136: data_o = 32'h00000000 /* 0x3100 */;
                3137: data_o = 32'h00000000 /* 0x3104 */;
                3138: data_o = 32'h00000000 /* 0x3108 */;
                3139: data_o = 32'h00000000 /* 0x310c */;
                3140: data_o = 32'h00000000 /* 0x3110 */;
                3141: data_o = 32'h00000000 /* 0x3114 */;
                3142: data_o = 32'h00000000 /* 0x3118 */;
                3143: data_o = 32'h00000000 /* 0x311c */;
                3144: data_o = 32'h00000000 /* 0x3120 */;
                3145: data_o = 32'h00000000 /* 0x3124 */;
                3146: data_o = 32'h00000000 /* 0x3128 */;
                3147: data_o = 32'h00000000 /* 0x312c */;
                3148: data_o = 32'h00000000 /* 0x3130 */;
                3149: data_o = 32'h00000000 /* 0x3134 */;
                3150: data_o = 32'h00000000 /* 0x3138 */;
                3151: data_o = 32'h00000000 /* 0x313c */;
                3152: data_o = 32'h00000000 /* 0x3140 */;
                3153: data_o = 32'h00000000 /* 0x3144 */;
                3154: data_o = 32'h00000000 /* 0x3148 */;
                3155: data_o = 32'h00000000 /* 0x314c */;
                3156: data_o = 32'h00000000 /* 0x3150 */;
                3157: data_o = 32'h00000000 /* 0x3154 */;
                3158: data_o = 32'h00000000 /* 0x3158 */;
                3159: data_o = 32'h00000000 /* 0x315c */;
                3160: data_o = 32'h00000000 /* 0x3160 */;
                3161: data_o = 32'h00000000 /* 0x3164 */;
                3162: data_o = 32'h00000000 /* 0x3168 */;
                3163: data_o = 32'h00000000 /* 0x316c */;
                3164: data_o = 32'h00000000 /* 0x3170 */;
                3165: data_o = 32'h00000000 /* 0x3174 */;
                3166: data_o = 32'h00000000 /* 0x3178 */;
                3167: data_o = 32'h00000000 /* 0x317c */;
                3168: data_o = 32'h00000000 /* 0x3180 */;
                3169: data_o = 32'h00000000 /* 0x3184 */;
                3170: data_o = 32'h00000000 /* 0x3188 */;
                3171: data_o = 32'h00000000 /* 0x318c */;
                3172: data_o = 32'h00000000 /* 0x3190 */;
                3173: data_o = 32'h00000000 /* 0x3194 */;
                3174: data_o = 32'h00000000 /* 0x3198 */;
                3175: data_o = 32'h00000000 /* 0x319c */;
                3176: data_o = 32'h00000000 /* 0x31a0 */;
                3177: data_o = 32'h00000000 /* 0x31a4 */;
                3178: data_o = 32'h00000000 /* 0x31a8 */;
                3179: data_o = 32'h00000000 /* 0x31ac */;
                3180: data_o = 32'h00000000 /* 0x31b0 */;
                3181: data_o = 32'h00000000 /* 0x31b4 */;
                3182: data_o = 32'h00000000 /* 0x31b8 */;
                3183: data_o = 32'h00000000 /* 0x31bc */;
                3184: data_o = 32'h00000000 /* 0x31c0 */;
                3185: data_o = 32'h00000000 /* 0x31c4 */;
                3186: data_o = 32'h00000000 /* 0x31c8 */;
                3187: data_o = 32'h00000000 /* 0x31cc */;
                3188: data_o = 32'h00000000 /* 0x31d0 */;
                3189: data_o = 32'h00000000 /* 0x31d4 */;
                3190: data_o = 32'h00000000 /* 0x31d8 */;
                3191: data_o = 32'h00000000 /* 0x31dc */;
                3192: data_o = 32'h00000000 /* 0x31e0 */;
                3193: data_o = 32'h00000000 /* 0x31e4 */;
                3194: data_o = 32'h00000000 /* 0x31e8 */;
                3195: data_o = 32'h00000000 /* 0x31ec */;
                3196: data_o = 32'h00000000 /* 0x31f0 */;
                3197: data_o = 32'h00000000 /* 0x31f4 */;
                3198: data_o = 32'h00000000 /* 0x31f8 */;
                3199: data_o = 32'h00000000 /* 0x31fc */;
                3200: data_o = 32'h00000000 /* 0x3200 */;
                3201: data_o = 32'h00000000 /* 0x3204 */;
                3202: data_o = 32'h00000000 /* 0x3208 */;
                3203: data_o = 32'h00000000 /* 0x320c */;
                3204: data_o = 32'h00000000 /* 0x3210 */;
                3205: data_o = 32'h00000000 /* 0x3214 */;
                3206: data_o = 32'h00000000 /* 0x3218 */;
                3207: data_o = 32'h00000000 /* 0x321c */;
                3208: data_o = 32'h00000000 /* 0x3220 */;
                3209: data_o = 32'h00000000 /* 0x3224 */;
                3210: data_o = 32'h00000000 /* 0x3228 */;
                3211: data_o = 32'h00000000 /* 0x322c */;
                3212: data_o = 32'h00000000 /* 0x3230 */;
                3213: data_o = 32'h00000000 /* 0x3234 */;
                3214: data_o = 32'h00000000 /* 0x3238 */;
                3215: data_o = 32'h00000000 /* 0x323c */;
                3216: data_o = 32'h00000000 /* 0x3240 */;
                3217: data_o = 32'h00000000 /* 0x3244 */;
                3218: data_o = 32'h00000000 /* 0x3248 */;
                3219: data_o = 32'h00000000 /* 0x324c */;
                3220: data_o = 32'h00000000 /* 0x3250 */;
                3221: data_o = 32'h00000000 /* 0x3254 */;
                3222: data_o = 32'h00000000 /* 0x3258 */;
                3223: data_o = 32'h00000000 /* 0x325c */;
                3224: data_o = 32'h00000000 /* 0x3260 */;
                3225: data_o = 32'h00000000 /* 0x3264 */;
                3226: data_o = 32'h00000000 /* 0x3268 */;
                3227: data_o = 32'h00000000 /* 0x326c */;
                3228: data_o = 32'h00000000 /* 0x3270 */;
                3229: data_o = 32'h00000000 /* 0x3274 */;
                3230: data_o = 32'h00000000 /* 0x3278 */;
                3231: data_o = 32'h00000000 /* 0x327c */;
                3232: data_o = 32'h00000000 /* 0x3280 */;
                3233: data_o = 32'h00000000 /* 0x3284 */;
                3234: data_o = 32'h00000000 /* 0x3288 */;
                3235: data_o = 32'h00000000 /* 0x328c */;
                3236: data_o = 32'h00000000 /* 0x3290 */;
                3237: data_o = 32'h00000000 /* 0x3294 */;
                3238: data_o = 32'h00000000 /* 0x3298 */;
                3239: data_o = 32'h00000000 /* 0x329c */;
                3240: data_o = 32'h00000000 /* 0x32a0 */;
                3241: data_o = 32'h00000000 /* 0x32a4 */;
                3242: data_o = 32'h00000000 /* 0x32a8 */;
                3243: data_o = 32'h00000000 /* 0x32ac */;
                3244: data_o = 32'h00000000 /* 0x32b0 */;
                3245: data_o = 32'h00000000 /* 0x32b4 */;
                3246: data_o = 32'h00000000 /* 0x32b8 */;
                3247: data_o = 32'h00000000 /* 0x32bc */;
                3248: data_o = 32'h00000000 /* 0x32c0 */;
                3249: data_o = 32'h00000000 /* 0x32c4 */;
                3250: data_o = 32'h00000000 /* 0x32c8 */;
                3251: data_o = 32'h00000000 /* 0x32cc */;
                3252: data_o = 32'h00000000 /* 0x32d0 */;
                3253: data_o = 32'h00000000 /* 0x32d4 */;
                3254: data_o = 32'h00000000 /* 0x32d8 */;
                3255: data_o = 32'h00000000 /* 0x32dc */;
                3256: data_o = 32'h00000000 /* 0x32e0 */;
                3257: data_o = 32'h00000000 /* 0x32e4 */;
                3258: data_o = 32'h00000000 /* 0x32e8 */;
                3259: data_o = 32'h00000000 /* 0x32ec */;
                3260: data_o = 32'h00000000 /* 0x32f0 */;
                3261: data_o = 32'h00000000 /* 0x32f4 */;
                3262: data_o = 32'h00000000 /* 0x32f8 */;
                3263: data_o = 32'h00000000 /* 0x32fc */;
                3264: data_o = 32'h00000000 /* 0x3300 */;
                3265: data_o = 32'h00000000 /* 0x3304 */;
                3266: data_o = 32'h00000000 /* 0x3308 */;
                3267: data_o = 32'h00000000 /* 0x330c */;
                3268: data_o = 32'h00000000 /* 0x3310 */;
                3269: data_o = 32'h00000000 /* 0x3314 */;
                3270: data_o = 32'h00000000 /* 0x3318 */;
                3271: data_o = 32'h00000000 /* 0x331c */;
                3272: data_o = 32'h00000000 /* 0x3320 */;
                3273: data_o = 32'h00000000 /* 0x3324 */;
                3274: data_o = 32'h00000000 /* 0x3328 */;
                3275: data_o = 32'h00000000 /* 0x332c */;
                3276: data_o = 32'h00000000 /* 0x3330 */;
                3277: data_o = 32'h00000000 /* 0x3334 */;
                3278: data_o = 32'h00000000 /* 0x3338 */;
                3279: data_o = 32'h00000000 /* 0x333c */;
                3280: data_o = 32'h00000000 /* 0x3340 */;
                3281: data_o = 32'h00000000 /* 0x3344 */;
                3282: data_o = 32'h00000000 /* 0x3348 */;
                3283: data_o = 32'h00000000 /* 0x334c */;
                3284: data_o = 32'h00000000 /* 0x3350 */;
                3285: data_o = 32'h00000000 /* 0x3354 */;
                3286: data_o = 32'h00000000 /* 0x3358 */;
                3287: data_o = 32'h00000000 /* 0x335c */;
                3288: data_o = 32'h00000000 /* 0x3360 */;
                3289: data_o = 32'h00000000 /* 0x3364 */;
                3290: data_o = 32'h00000000 /* 0x3368 */;
                3291: data_o = 32'h00000000 /* 0x336c */;
                3292: data_o = 32'h00000000 /* 0x3370 */;
                3293: data_o = 32'h00000000 /* 0x3374 */;
                3294: data_o = 32'h00000000 /* 0x3378 */;
                3295: data_o = 32'h00000000 /* 0x337c */;
                3296: data_o = 32'h00000000 /* 0x3380 */;
                3297: data_o = 32'h00000000 /* 0x3384 */;
                3298: data_o = 32'h00000000 /* 0x3388 */;
                3299: data_o = 32'h00000000 /* 0x338c */;
                3300: data_o = 32'h00000000 /* 0x3390 */;
                3301: data_o = 32'h00000000 /* 0x3394 */;
                3302: data_o = 32'h00000000 /* 0x3398 */;
                3303: data_o = 32'h00000000 /* 0x339c */;
                3304: data_o = 32'h00000000 /* 0x33a0 */;
                3305: data_o = 32'h00000000 /* 0x33a4 */;
                3306: data_o = 32'h00000000 /* 0x33a8 */;
                3307: data_o = 32'h00000000 /* 0x33ac */;
                3308: data_o = 32'h00000000 /* 0x33b0 */;
                3309: data_o = 32'h00000000 /* 0x33b4 */;
                3310: data_o = 32'h00000000 /* 0x33b8 */;
                3311: data_o = 32'h00000000 /* 0x33bc */;
                3312: data_o = 32'h00000000 /* 0x33c0 */;
                3313: data_o = 32'h00000000 /* 0x33c4 */;
                3314: data_o = 32'h00000000 /* 0x33c8 */;
                3315: data_o = 32'h00000000 /* 0x33cc */;
                3316: data_o = 32'h00000000 /* 0x33d0 */;
                3317: data_o = 32'h00000000 /* 0x33d4 */;
                3318: data_o = 32'h00000000 /* 0x33d8 */;
                3319: data_o = 32'h00000000 /* 0x33dc */;
                3320: data_o = 32'h00000000 /* 0x33e0 */;
                3321: data_o = 32'h00000000 /* 0x33e4 */;
                3322: data_o = 32'h00000000 /* 0x33e8 */;
                3323: data_o = 32'h00000000 /* 0x33ec */;
                3324: data_o = 32'h00000000 /* 0x33f0 */;
                3325: data_o = 32'h00000000 /* 0x33f4 */;
                3326: data_o = 32'h00000000 /* 0x33f8 */;
                3327: data_o = 32'h00000000 /* 0x33fc */;
                3328: data_o = 32'h00000000 /* 0x3400 */;
                3329: data_o = 32'h00000000 /* 0x3404 */;
                3330: data_o = 32'h00000000 /* 0x3408 */;
                3331: data_o = 32'h00000000 /* 0x340c */;
                3332: data_o = 32'h00000000 /* 0x3410 */;
                3333: data_o = 32'h00000000 /* 0x3414 */;
                3334: data_o = 32'h00000000 /* 0x3418 */;
                3335: data_o = 32'h00000000 /* 0x341c */;
                3336: data_o = 32'h00000000 /* 0x3420 */;
                3337: data_o = 32'h00000000 /* 0x3424 */;
                3338: data_o = 32'h00000000 /* 0x3428 */;
                3339: data_o = 32'h00000000 /* 0x342c */;
                3340: data_o = 32'h00000000 /* 0x3430 */;
                3341: data_o = 32'h00000000 /* 0x3434 */;
                3342: data_o = 32'h00000000 /* 0x3438 */;
                3343: data_o = 32'h00000000 /* 0x343c */;
                3344: data_o = 32'h00000000 /* 0x3440 */;
                3345: data_o = 32'h00000000 /* 0x3444 */;
                3346: data_o = 32'h00000000 /* 0x3448 */;
                3347: data_o = 32'h00000000 /* 0x344c */;
                3348: data_o = 32'h00000000 /* 0x3450 */;
                3349: data_o = 32'h00000000 /* 0x3454 */;
                3350: data_o = 32'h00000000 /* 0x3458 */;
                3351: data_o = 32'h00000000 /* 0x345c */;
                3352: data_o = 32'h00000000 /* 0x3460 */;
                3353: data_o = 32'h00000000 /* 0x3464 */;
                3354: data_o = 32'h00000000 /* 0x3468 */;
                3355: data_o = 32'h00000000 /* 0x346c */;
                3356: data_o = 32'h00000000 /* 0x3470 */;
                3357: data_o = 32'h00000000 /* 0x3474 */;
                3358: data_o = 32'h00000000 /* 0x3478 */;
                3359: data_o = 32'h00000000 /* 0x347c */;
                3360: data_o = 32'h00000000 /* 0x3480 */;
                3361: data_o = 32'h00000000 /* 0x3484 */;
                3362: data_o = 32'h00000000 /* 0x3488 */;
                3363: data_o = 32'h00000000 /* 0x348c */;
                3364: data_o = 32'h00000000 /* 0x3490 */;
                3365: data_o = 32'h00000000 /* 0x3494 */;
                3366: data_o = 32'h00000000 /* 0x3498 */;
                3367: data_o = 32'h00000000 /* 0x349c */;
                3368: data_o = 32'h00000000 /* 0x34a0 */;
                3369: data_o = 32'h00000000 /* 0x34a4 */;
                3370: data_o = 32'h00000000 /* 0x34a8 */;
                3371: data_o = 32'h00000000 /* 0x34ac */;
                3372: data_o = 32'h00000000 /* 0x34b0 */;
                3373: data_o = 32'h00000000 /* 0x34b4 */;
                3374: data_o = 32'h00000000 /* 0x34b8 */;
                3375: data_o = 32'h00000000 /* 0x34bc */;
                3376: data_o = 32'h00000000 /* 0x34c0 */;
                3377: data_o = 32'h00000000 /* 0x34c4 */;
                3378: data_o = 32'h00000000 /* 0x34c8 */;
                3379: data_o = 32'h00000000 /* 0x34cc */;
                3380: data_o = 32'h00000000 /* 0x34d0 */;
                3381: data_o = 32'h00000000 /* 0x34d4 */;
                3382: data_o = 32'h00000000 /* 0x34d8 */;
                3383: data_o = 32'h00000000 /* 0x34dc */;
                3384: data_o = 32'h00000000 /* 0x34e0 */;
                3385: data_o = 32'h00000000 /* 0x34e4 */;
                3386: data_o = 32'h00000000 /* 0x34e8 */;
                3387: data_o = 32'h00000000 /* 0x34ec */;
                3388: data_o = 32'h00000000 /* 0x34f0 */;
                3389: data_o = 32'h00000000 /* 0x34f4 */;
                3390: data_o = 32'h00000000 /* 0x34f8 */;
                3391: data_o = 32'h00000000 /* 0x34fc */;
                3392: data_o = 32'h00000000 /* 0x3500 */;
                3393: data_o = 32'h00000000 /* 0x3504 */;
                3394: data_o = 32'h00000000 /* 0x3508 */;
                3395: data_o = 32'h00000000 /* 0x350c */;
                3396: data_o = 32'h00000000 /* 0x3510 */;
                3397: data_o = 32'h00000000 /* 0x3514 */;
                3398: data_o = 32'h00000000 /* 0x3518 */;
                3399: data_o = 32'h00000000 /* 0x351c */;
                3400: data_o = 32'h00000000 /* 0x3520 */;
                3401: data_o = 32'h00000000 /* 0x3524 */;
                3402: data_o = 32'h00000000 /* 0x3528 */;
                3403: data_o = 32'h00000000 /* 0x352c */;
                3404: data_o = 32'h00000000 /* 0x3530 */;
                3405: data_o = 32'h00000000 /* 0x3534 */;
                3406: data_o = 32'h00000000 /* 0x3538 */;
                3407: data_o = 32'h00000000 /* 0x353c */;
                3408: data_o = 32'h00000000 /* 0x3540 */;
                3409: data_o = 32'h00000000 /* 0x3544 */;
                3410: data_o = 32'h00000000 /* 0x3548 */;
                3411: data_o = 32'h00000000 /* 0x354c */;
                3412: data_o = 32'h00000000 /* 0x3550 */;
                3413: data_o = 32'h00000000 /* 0x3554 */;
                3414: data_o = 32'h00000000 /* 0x3558 */;
                3415: data_o = 32'h00000000 /* 0x355c */;
                3416: data_o = 32'h00000000 /* 0x3560 */;
                3417: data_o = 32'h00000000 /* 0x3564 */;
                3418: data_o = 32'h00000000 /* 0x3568 */;
                3419: data_o = 32'h00000000 /* 0x356c */;
                3420: data_o = 32'h00000000 /* 0x3570 */;
                3421: data_o = 32'h00000000 /* 0x3574 */;
                3422: data_o = 32'h00000000 /* 0x3578 */;
                3423: data_o = 32'h00000000 /* 0x357c */;
                3424: data_o = 32'h00000000 /* 0x3580 */;
                3425: data_o = 32'h00000000 /* 0x3584 */;
                3426: data_o = 32'h00000000 /* 0x3588 */;
                3427: data_o = 32'h00000000 /* 0x358c */;
                3428: data_o = 32'h00000000 /* 0x3590 */;
                3429: data_o = 32'h00000000 /* 0x3594 */;
                3430: data_o = 32'h00000000 /* 0x3598 */;
                3431: data_o = 32'h00000000 /* 0x359c */;
                3432: data_o = 32'h00000000 /* 0x35a0 */;
                3433: data_o = 32'h00000000 /* 0x35a4 */;
                3434: data_o = 32'h00000000 /* 0x35a8 */;
                3435: data_o = 32'h00000000 /* 0x35ac */;
                3436: data_o = 32'h00000000 /* 0x35b0 */;
                3437: data_o = 32'h00000000 /* 0x35b4 */;
                3438: data_o = 32'h00000000 /* 0x35b8 */;
                3439: data_o = 32'h00000000 /* 0x35bc */;
                3440: data_o = 32'h00000000 /* 0x35c0 */;
                3441: data_o = 32'h00000000 /* 0x35c4 */;
                3442: data_o = 32'h00000000 /* 0x35c8 */;
                3443: data_o = 32'h00000000 /* 0x35cc */;
                3444: data_o = 32'h00000000 /* 0x35d0 */;
                3445: data_o = 32'h00000000 /* 0x35d4 */;
                3446: data_o = 32'h00000000 /* 0x35d8 */;
                3447: data_o = 32'h00000000 /* 0x35dc */;
                3448: data_o = 32'h00000000 /* 0x35e0 */;
                3449: data_o = 32'h00000000 /* 0x35e4 */;
                3450: data_o = 32'h00000000 /* 0x35e8 */;
                3451: data_o = 32'h00000000 /* 0x35ec */;
                3452: data_o = 32'h00000000 /* 0x35f0 */;
                3453: data_o = 32'h00000000 /* 0x35f4 */;
                3454: data_o = 32'h00000000 /* 0x35f8 */;
                3455: data_o = 32'h00000000 /* 0x35fc */;
                3456: data_o = 32'h00000000 /* 0x3600 */;
                3457: data_o = 32'h00000000 /* 0x3604 */;
                3458: data_o = 32'h00000000 /* 0x3608 */;
                3459: data_o = 32'h00000000 /* 0x360c */;
                3460: data_o = 32'h00000000 /* 0x3610 */;
                3461: data_o = 32'h00000000 /* 0x3614 */;
                3462: data_o = 32'h00000000 /* 0x3618 */;
                3463: data_o = 32'h00000000 /* 0x361c */;
                3464: data_o = 32'h00000000 /* 0x3620 */;
                3465: data_o = 32'h00000000 /* 0x3624 */;
                3466: data_o = 32'h00000000 /* 0x3628 */;
                3467: data_o = 32'h00000000 /* 0x362c */;
                3468: data_o = 32'h00000000 /* 0x3630 */;
                3469: data_o = 32'h00000000 /* 0x3634 */;
                3470: data_o = 32'h00000000 /* 0x3638 */;
                3471: data_o = 32'h00000000 /* 0x363c */;
                3472: data_o = 32'h00000000 /* 0x3640 */;
                3473: data_o = 32'h00000000 /* 0x3644 */;
                3474: data_o = 32'h00000000 /* 0x3648 */;
                3475: data_o = 32'h00000000 /* 0x364c */;
                3476: data_o = 32'h00000000 /* 0x3650 */;
                3477: data_o = 32'h00000000 /* 0x3654 */;
                3478: data_o = 32'h00000000 /* 0x3658 */;
                3479: data_o = 32'h00000000 /* 0x365c */;
                3480: data_o = 32'h00000000 /* 0x3660 */;
                3481: data_o = 32'h00000000 /* 0x3664 */;
                3482: data_o = 32'h00000000 /* 0x3668 */;
                3483: data_o = 32'h00000000 /* 0x366c */;
                3484: data_o = 32'h00000000 /* 0x3670 */;
                3485: data_o = 32'h00000000 /* 0x3674 */;
                3486: data_o = 32'h00000000 /* 0x3678 */;
                3487: data_o = 32'h00000000 /* 0x367c */;
                3488: data_o = 32'h00000000 /* 0x3680 */;
                3489: data_o = 32'h00000000 /* 0x3684 */;
                3490: data_o = 32'h00000000 /* 0x3688 */;
                3491: data_o = 32'h00000000 /* 0x368c */;
                3492: data_o = 32'h00000000 /* 0x3690 */;
                3493: data_o = 32'h00000000 /* 0x3694 */;
                3494: data_o = 32'h00000000 /* 0x3698 */;
                3495: data_o = 32'h00000000 /* 0x369c */;
                3496: data_o = 32'h00000000 /* 0x36a0 */;
                3497: data_o = 32'h00000000 /* 0x36a4 */;
                3498: data_o = 32'h00000000 /* 0x36a8 */;
                3499: data_o = 32'h00000000 /* 0x36ac */;
                3500: data_o = 32'h00000000 /* 0x36b0 */;
                3501: data_o = 32'h00000000 /* 0x36b4 */;
                3502: data_o = 32'h00000000 /* 0x36b8 */;
                3503: data_o = 32'h00000000 /* 0x36bc */;
                3504: data_o = 32'h00000000 /* 0x36c0 */;
                3505: data_o = 32'h00000000 /* 0x36c4 */;
                3506: data_o = 32'h00000000 /* 0x36c8 */;
                3507: data_o = 32'h00000000 /* 0x36cc */;
                3508: data_o = 32'h00000000 /* 0x36d0 */;
                3509: data_o = 32'h00000000 /* 0x36d4 */;
                3510: data_o = 32'h00000000 /* 0x36d8 */;
                3511: data_o = 32'h00000000 /* 0x36dc */;
                3512: data_o = 32'h00000000 /* 0x36e0 */;
                3513: data_o = 32'h00000000 /* 0x36e4 */;
                3514: data_o = 32'h00000000 /* 0x36e8 */;
                3515: data_o = 32'h00000000 /* 0x36ec */;
                3516: data_o = 32'h00000000 /* 0x36f0 */;
                3517: data_o = 32'h00000000 /* 0x36f4 */;
                3518: data_o = 32'h00000000 /* 0x36f8 */;
                3519: data_o = 32'h00000000 /* 0x36fc */;
                3520: data_o = 32'h00000000 /* 0x3700 */;
                3521: data_o = 32'h00000000 /* 0x3704 */;
                3522: data_o = 32'h00000000 /* 0x3708 */;
                3523: data_o = 32'h00000000 /* 0x370c */;
                3524: data_o = 32'h00000000 /* 0x3710 */;
                3525: data_o = 32'h00000000 /* 0x3714 */;
                3526: data_o = 32'h00000000 /* 0x3718 */;
                3527: data_o = 32'h00000000 /* 0x371c */;
                3528: data_o = 32'h00000000 /* 0x3720 */;
                3529: data_o = 32'h00000000 /* 0x3724 */;
                3530: data_o = 32'h00000000 /* 0x3728 */;
                3531: data_o = 32'h00000000 /* 0x372c */;
                3532: data_o = 32'h00000000 /* 0x3730 */;
                3533: data_o = 32'h00000000 /* 0x3734 */;
                3534: data_o = 32'h00000000 /* 0x3738 */;
                3535: data_o = 32'h00000000 /* 0x373c */;
                3536: data_o = 32'h00000000 /* 0x3740 */;
                3537: data_o = 32'h00000000 /* 0x3744 */;
                3538: data_o = 32'h00000000 /* 0x3748 */;
                3539: data_o = 32'h00000000 /* 0x374c */;
                3540: data_o = 32'h00000000 /* 0x3750 */;
                3541: data_o = 32'h00000000 /* 0x3754 */;
                3542: data_o = 32'h00000000 /* 0x3758 */;
                3543: data_o = 32'h00000000 /* 0x375c */;
                3544: data_o = 32'h00000000 /* 0x3760 */;
                3545: data_o = 32'h00000000 /* 0x3764 */;
                3546: data_o = 32'h00000000 /* 0x3768 */;
                3547: data_o = 32'h00000000 /* 0x376c */;
                3548: data_o = 32'h00000000 /* 0x3770 */;
                3549: data_o = 32'h00000000 /* 0x3774 */;
                3550: data_o = 32'h00000000 /* 0x3778 */;
                3551: data_o = 32'h00000000 /* 0x377c */;
                3552: data_o = 32'h00000000 /* 0x3780 */;
                3553: data_o = 32'h00000000 /* 0x3784 */;
                3554: data_o = 32'h00000000 /* 0x3788 */;
                3555: data_o = 32'h00000000 /* 0x378c */;
                3556: data_o = 32'h00000000 /* 0x3790 */;
                3557: data_o = 32'h00000000 /* 0x3794 */;
                3558: data_o = 32'h00000000 /* 0x3798 */;
                3559: data_o = 32'h00000000 /* 0x379c */;
                3560: data_o = 32'h00000000 /* 0x37a0 */;
                3561: data_o = 32'h00000000 /* 0x37a4 */;
                3562: data_o = 32'h00000000 /* 0x37a8 */;
                3563: data_o = 32'h00000000 /* 0x37ac */;
                3564: data_o = 32'h00000000 /* 0x37b0 */;
                3565: data_o = 32'h00000000 /* 0x37b4 */;
                3566: data_o = 32'h00000000 /* 0x37b8 */;
                3567: data_o = 32'h00000000 /* 0x37bc */;
                3568: data_o = 32'h00000000 /* 0x37c0 */;
                3569: data_o = 32'h00000000 /* 0x37c4 */;
                3570: data_o = 32'h00000000 /* 0x37c8 */;
                3571: data_o = 32'h00000000 /* 0x37cc */;
                3572: data_o = 32'h00000000 /* 0x37d0 */;
                3573: data_o = 32'h00000000 /* 0x37d4 */;
                3574: data_o = 32'h00000000 /* 0x37d8 */;
                3575: data_o = 32'h00000000 /* 0x37dc */;
                3576: data_o = 32'h00000000 /* 0x37e0 */;
                3577: data_o = 32'h00000000 /* 0x37e4 */;
                3578: data_o = 32'h00000000 /* 0x37e8 */;
                3579: data_o = 32'h00000000 /* 0x37ec */;
                3580: data_o = 32'h00000000 /* 0x37f0 */;
                3581: data_o = 32'h00000000 /* 0x37f4 */;
                3582: data_o = 32'h00000000 /* 0x37f8 */;
                3583: data_o = 32'h00000000 /* 0x37fc */;
                3584: data_o = 32'h00000000 /* 0x3800 */;
                3585: data_o = 32'h00000000 /* 0x3804 */;
                3586: data_o = 32'h00000000 /* 0x3808 */;
                3587: data_o = 32'h00000000 /* 0x380c */;
                3588: data_o = 32'h00000000 /* 0x3810 */;
                3589: data_o = 32'h00000000 /* 0x3814 */;
                3590: data_o = 32'h00000000 /* 0x3818 */;
                3591: data_o = 32'h00000000 /* 0x381c */;
                3592: data_o = 32'h00000000 /* 0x3820 */;
                3593: data_o = 32'h00000000 /* 0x3824 */;
                3594: data_o = 32'h00000000 /* 0x3828 */;
                3595: data_o = 32'h00000000 /* 0x382c */;
                3596: data_o = 32'h00000000 /* 0x3830 */;
                3597: data_o = 32'h00000000 /* 0x3834 */;
                3598: data_o = 32'h00000000 /* 0x3838 */;
                3599: data_o = 32'h00000000 /* 0x383c */;
                3600: data_o = 32'h00000000 /* 0x3840 */;
                3601: data_o = 32'h00000000 /* 0x3844 */;
                3602: data_o = 32'h00000000 /* 0x3848 */;
                3603: data_o = 32'h00000000 /* 0x384c */;
                3604: data_o = 32'h00000000 /* 0x3850 */;
                3605: data_o = 32'h00000000 /* 0x3854 */;
                3606: data_o = 32'h00000000 /* 0x3858 */;
                3607: data_o = 32'h00000000 /* 0x385c */;
                3608: data_o = 32'h00000000 /* 0x3860 */;
                3609: data_o = 32'h00000000 /* 0x3864 */;
                3610: data_o = 32'h00000000 /* 0x3868 */;
                3611: data_o = 32'h00000000 /* 0x386c */;
                3612: data_o = 32'h00000000 /* 0x3870 */;
                3613: data_o = 32'h00000000 /* 0x3874 */;
                3614: data_o = 32'h00000000 /* 0x3878 */;
                3615: data_o = 32'h00000000 /* 0x387c */;
                3616: data_o = 32'h00000000 /* 0x3880 */;
                3617: data_o = 32'h00000000 /* 0x3884 */;
                3618: data_o = 32'h00000000 /* 0x3888 */;
                3619: data_o = 32'h00000000 /* 0x388c */;
                3620: data_o = 32'h00000000 /* 0x3890 */;
                3621: data_o = 32'h00000000 /* 0x3894 */;
                3622: data_o = 32'h00000000 /* 0x3898 */;
                3623: data_o = 32'h00000000 /* 0x389c */;
                3624: data_o = 32'h00000000 /* 0x38a0 */;
                3625: data_o = 32'h00000000 /* 0x38a4 */;
                3626: data_o = 32'h00000000 /* 0x38a8 */;
                3627: data_o = 32'h00000000 /* 0x38ac */;
                3628: data_o = 32'h00000000 /* 0x38b0 */;
                3629: data_o = 32'h00000000 /* 0x38b4 */;
                3630: data_o = 32'h00000000 /* 0x38b8 */;
                3631: data_o = 32'h00000000 /* 0x38bc */;
                3632: data_o = 32'h00000000 /* 0x38c0 */;
                3633: data_o = 32'h00000000 /* 0x38c4 */;
                3634: data_o = 32'h00000000 /* 0x38c8 */;
                3635: data_o = 32'h00000000 /* 0x38cc */;
                3636: data_o = 32'h00000000 /* 0x38d0 */;
                3637: data_o = 32'h00000000 /* 0x38d4 */;
                3638: data_o = 32'h00000000 /* 0x38d8 */;
                3639: data_o = 32'h00000000 /* 0x38dc */;
                3640: data_o = 32'h00000000 /* 0x38e0 */;
                3641: data_o = 32'h00000000 /* 0x38e4 */;
                3642: data_o = 32'h00000000 /* 0x38e8 */;
                3643: data_o = 32'h00000000 /* 0x38ec */;
                3644: data_o = 32'h00000000 /* 0x38f0 */;
                3645: data_o = 32'h00000000 /* 0x38f4 */;
                3646: data_o = 32'h00000000 /* 0x38f8 */;
                3647: data_o = 32'h00000000 /* 0x38fc */;
                3648: data_o = 32'h00000000 /* 0x3900 */;
                3649: data_o = 32'h00000000 /* 0x3904 */;
                3650: data_o = 32'h00000000 /* 0x3908 */;
                3651: data_o = 32'h00000000 /* 0x390c */;
                3652: data_o = 32'h00000000 /* 0x3910 */;
                3653: data_o = 32'h00000000 /* 0x3914 */;
                3654: data_o = 32'h00000000 /* 0x3918 */;
                3655: data_o = 32'h00000000 /* 0x391c */;
                3656: data_o = 32'h00000000 /* 0x3920 */;
                3657: data_o = 32'h00000000 /* 0x3924 */;
                3658: data_o = 32'h00000000 /* 0x3928 */;
                3659: data_o = 32'h00000000 /* 0x392c */;
                3660: data_o = 32'h00000000 /* 0x3930 */;
                3661: data_o = 32'h00000000 /* 0x3934 */;
                3662: data_o = 32'h00000000 /* 0x3938 */;
                3663: data_o = 32'h00000000 /* 0x393c */;
                3664: data_o = 32'h00000000 /* 0x3940 */;
                3665: data_o = 32'h00000000 /* 0x3944 */;
                3666: data_o = 32'h00000000 /* 0x3948 */;
                3667: data_o = 32'h00000000 /* 0x394c */;
                3668: data_o = 32'h00000000 /* 0x3950 */;
                3669: data_o = 32'h00000000 /* 0x3954 */;
                3670: data_o = 32'h00000000 /* 0x3958 */;
                3671: data_o = 32'h00000000 /* 0x395c */;
                3672: data_o = 32'h00000000 /* 0x3960 */;
                3673: data_o = 32'h00000000 /* 0x3964 */;
                3674: data_o = 32'h00000000 /* 0x3968 */;
                3675: data_o = 32'h00000000 /* 0x396c */;
                3676: data_o = 32'h00000000 /* 0x3970 */;
                3677: data_o = 32'h00000000 /* 0x3974 */;
                3678: data_o = 32'h00000000 /* 0x3978 */;
                3679: data_o = 32'h00000000 /* 0x397c */;
                3680: data_o = 32'h00000000 /* 0x3980 */;
                3681: data_o = 32'h00000000 /* 0x3984 */;
                3682: data_o = 32'h00000000 /* 0x3988 */;
                3683: data_o = 32'h00000000 /* 0x398c */;
                3684: data_o = 32'h00000000 /* 0x3990 */;
                3685: data_o = 32'h00000000 /* 0x3994 */;
                3686: data_o = 32'h00000000 /* 0x3998 */;
                3687: data_o = 32'h00000000 /* 0x399c */;
                3688: data_o = 32'h00000000 /* 0x39a0 */;
                3689: data_o = 32'h00000000 /* 0x39a4 */;
                3690: data_o = 32'h00000000 /* 0x39a8 */;
                3691: data_o = 32'h00000000 /* 0x39ac */;
                3692: data_o = 32'h00000000 /* 0x39b0 */;
                3693: data_o = 32'h00000000 /* 0x39b4 */;
                3694: data_o = 32'h00000000 /* 0x39b8 */;
                3695: data_o = 32'h00000000 /* 0x39bc */;
                3696: data_o = 32'h00000000 /* 0x39c0 */;
                3697: data_o = 32'h00000000 /* 0x39c4 */;
                3698: data_o = 32'h00000000 /* 0x39c8 */;
                3699: data_o = 32'h00000000 /* 0x39cc */;
                3700: data_o = 32'h00000000 /* 0x39d0 */;
                3701: data_o = 32'h00000000 /* 0x39d4 */;
                3702: data_o = 32'h00000000 /* 0x39d8 */;
                3703: data_o = 32'h00000000 /* 0x39dc */;
                3704: data_o = 32'h00000000 /* 0x39e0 */;
                3705: data_o = 32'h00000000 /* 0x39e4 */;
                3706: data_o = 32'h00000000 /* 0x39e8 */;
                3707: data_o = 32'h00000000 /* 0x39ec */;
                3708: data_o = 32'h00000000 /* 0x39f0 */;
                3709: data_o = 32'h00000000 /* 0x39f4 */;
                3710: data_o = 32'h00000000 /* 0x39f8 */;
                3711: data_o = 32'h00000000 /* 0x39fc */;
                3712: data_o = 32'h00000000 /* 0x3a00 */;
                3713: data_o = 32'h00000000 /* 0x3a04 */;
                3714: data_o = 32'h00000000 /* 0x3a08 */;
                3715: data_o = 32'h00000000 /* 0x3a0c */;
                3716: data_o = 32'h00000000 /* 0x3a10 */;
                3717: data_o = 32'h00000000 /* 0x3a14 */;
                3718: data_o = 32'h00000000 /* 0x3a18 */;
                3719: data_o = 32'h00000000 /* 0x3a1c */;
                3720: data_o = 32'h00000000 /* 0x3a20 */;
                3721: data_o = 32'h00000000 /* 0x3a24 */;
                3722: data_o = 32'h00000000 /* 0x3a28 */;
                3723: data_o = 32'h00000000 /* 0x3a2c */;
                3724: data_o = 32'h00000000 /* 0x3a30 */;
                3725: data_o = 32'h00000000 /* 0x3a34 */;
                3726: data_o = 32'h00000000 /* 0x3a38 */;
                3727: data_o = 32'h00000000 /* 0x3a3c */;
                3728: data_o = 32'h00000000 /* 0x3a40 */;
                3729: data_o = 32'h00000000 /* 0x3a44 */;
                3730: data_o = 32'h00000000 /* 0x3a48 */;
                3731: data_o = 32'h00000000 /* 0x3a4c */;
                3732: data_o = 32'h00000000 /* 0x3a50 */;
                3733: data_o = 32'h00000000 /* 0x3a54 */;
                3734: data_o = 32'h00000000 /* 0x3a58 */;
                3735: data_o = 32'h00000000 /* 0x3a5c */;
                3736: data_o = 32'h00000000 /* 0x3a60 */;
                3737: data_o = 32'h00000000 /* 0x3a64 */;
                3738: data_o = 32'h00000000 /* 0x3a68 */;
                3739: data_o = 32'h00000000 /* 0x3a6c */;
                3740: data_o = 32'h00000000 /* 0x3a70 */;
                3741: data_o = 32'h00000000 /* 0x3a74 */;
                3742: data_o = 32'h00000000 /* 0x3a78 */;
                3743: data_o = 32'h00000000 /* 0x3a7c */;
                3744: data_o = 32'h00000000 /* 0x3a80 */;
                3745: data_o = 32'h00000000 /* 0x3a84 */;
                3746: data_o = 32'h00000000 /* 0x3a88 */;
                3747: data_o = 32'h00000000 /* 0x3a8c */;
                3748: data_o = 32'h00000000 /* 0x3a90 */;
                3749: data_o = 32'h00000000 /* 0x3a94 */;
                3750: data_o = 32'h00000000 /* 0x3a98 */;
                3751: data_o = 32'h00000000 /* 0x3a9c */;
                3752: data_o = 32'h00000000 /* 0x3aa0 */;
                3753: data_o = 32'h00000000 /* 0x3aa4 */;
                3754: data_o = 32'h00000000 /* 0x3aa8 */;
                3755: data_o = 32'h00000000 /* 0x3aac */;
                3756: data_o = 32'h00000000 /* 0x3ab0 */;
                3757: data_o = 32'h00000000 /* 0x3ab4 */;
                3758: data_o = 32'h00000000 /* 0x3ab8 */;
                3759: data_o = 32'h00000000 /* 0x3abc */;
                3760: data_o = 32'h00000000 /* 0x3ac0 */;
                3761: data_o = 32'h00000000 /* 0x3ac4 */;
                3762: data_o = 32'h00000000 /* 0x3ac8 */;
                3763: data_o = 32'h00000000 /* 0x3acc */;
                3764: data_o = 32'h00000000 /* 0x3ad0 */;
                3765: data_o = 32'h00000000 /* 0x3ad4 */;
                3766: data_o = 32'h00000000 /* 0x3ad8 */;
                3767: data_o = 32'h00000000 /* 0x3adc */;
                3768: data_o = 32'h00000000 /* 0x3ae0 */;
                3769: data_o = 32'h00000000 /* 0x3ae4 */;
                3770: data_o = 32'h00000000 /* 0x3ae8 */;
                3771: data_o = 32'h00000000 /* 0x3aec */;
                3772: data_o = 32'h00000000 /* 0x3af0 */;
                3773: data_o = 32'h00000000 /* 0x3af4 */;
                3774: data_o = 32'h00000000 /* 0x3af8 */;
                3775: data_o = 32'h00000000 /* 0x3afc */;
                3776: data_o = 32'h00000000 /* 0x3b00 */;
                3777: data_o = 32'h00000000 /* 0x3b04 */;
                3778: data_o = 32'h00000000 /* 0x3b08 */;
                3779: data_o = 32'h00000000 /* 0x3b0c */;
                3780: data_o = 32'h00000000 /* 0x3b10 */;
                3781: data_o = 32'h00000000 /* 0x3b14 */;
                3782: data_o = 32'h00000000 /* 0x3b18 */;
                3783: data_o = 32'h00000000 /* 0x3b1c */;
                3784: data_o = 32'h00000000 /* 0x3b20 */;
                3785: data_o = 32'h00000000 /* 0x3b24 */;
                3786: data_o = 32'h00000000 /* 0x3b28 */;
                3787: data_o = 32'h00000000 /* 0x3b2c */;
                3788: data_o = 32'h00000000 /* 0x3b30 */;
                3789: data_o = 32'h00000000 /* 0x3b34 */;
                3790: data_o = 32'h00000000 /* 0x3b38 */;
                3791: data_o = 32'h00000000 /* 0x3b3c */;
                3792: data_o = 32'h00000000 /* 0x3b40 */;
                3793: data_o = 32'h00000000 /* 0x3b44 */;
                3794: data_o = 32'h00000000 /* 0x3b48 */;
                3795: data_o = 32'h00000000 /* 0x3b4c */;
                3796: data_o = 32'h00000000 /* 0x3b50 */;
                3797: data_o = 32'h00000000 /* 0x3b54 */;
                3798: data_o = 32'h00000000 /* 0x3b58 */;
                3799: data_o = 32'h00000000 /* 0x3b5c */;
                3800: data_o = 32'h00000000 /* 0x3b60 */;
                3801: data_o = 32'h00000000 /* 0x3b64 */;
                3802: data_o = 32'h00000000 /* 0x3b68 */;
                3803: data_o = 32'h00000000 /* 0x3b6c */;
                3804: data_o = 32'h00000000 /* 0x3b70 */;
                3805: data_o = 32'h00000000 /* 0x3b74 */;
                3806: data_o = 32'h00000000 /* 0x3b78 */;
                3807: data_o = 32'h00000000 /* 0x3b7c */;
                3808: data_o = 32'h00000000 /* 0x3b80 */;
                3809: data_o = 32'h00000000 /* 0x3b84 */;
                3810: data_o = 32'h00000000 /* 0x3b88 */;
                3811: data_o = 32'h00000000 /* 0x3b8c */;
                3812: data_o = 32'h00000000 /* 0x3b90 */;
                3813: data_o = 32'h00000000 /* 0x3b94 */;
                3814: data_o = 32'h00000000 /* 0x3b98 */;
                3815: data_o = 32'h00000000 /* 0x3b9c */;
                3816: data_o = 32'h00000000 /* 0x3ba0 */;
                3817: data_o = 32'h00000000 /* 0x3ba4 */;
                3818: data_o = 32'h00000000 /* 0x3ba8 */;
                3819: data_o = 32'h00000000 /* 0x3bac */;
                3820: data_o = 32'h00000000 /* 0x3bb0 */;
                3821: data_o = 32'h00000000 /* 0x3bb4 */;
                3822: data_o = 32'h00000000 /* 0x3bb8 */;
                3823: data_o = 32'h00000000 /* 0x3bbc */;
                3824: data_o = 32'h00000000 /* 0x3bc0 */;
                3825: data_o = 32'h00000000 /* 0x3bc4 */;
                3826: data_o = 32'h00000000 /* 0x3bc8 */;
                3827: data_o = 32'h00000000 /* 0x3bcc */;
                3828: data_o = 32'h00000000 /* 0x3bd0 */;
                3829: data_o = 32'h00000000 /* 0x3bd4 */;
                3830: data_o = 32'h00000000 /* 0x3bd8 */;
                3831: data_o = 32'h00000000 /* 0x3bdc */;
                3832: data_o = 32'h00000000 /* 0x3be0 */;
                3833: data_o = 32'h00000000 /* 0x3be4 */;
                3834: data_o = 32'h00000000 /* 0x3be8 */;
                3835: data_o = 32'h00000000 /* 0x3bec */;
                3836: data_o = 32'h00000000 /* 0x3bf0 */;
                3837: data_o = 32'h00000000 /* 0x3bf4 */;
                3838: data_o = 32'h00000000 /* 0x3bf8 */;
                3839: data_o = 32'h00000000 /* 0x3bfc */;
                3840: data_o = 32'h00000000 /* 0x3c00 */;
                3841: data_o = 32'h00000000 /* 0x3c04 */;
                3842: data_o = 32'h00000000 /* 0x3c08 */;
                3843: data_o = 32'h00000000 /* 0x3c0c */;
                3844: data_o = 32'h00000000 /* 0x3c10 */;
                3845: data_o = 32'h00000000 /* 0x3c14 */;
                3846: data_o = 32'h00000000 /* 0x3c18 */;
                3847: data_o = 32'h00000000 /* 0x3c1c */;
                3848: data_o = 32'h00000000 /* 0x3c20 */;
                3849: data_o = 32'h00000000 /* 0x3c24 */;
                3850: data_o = 32'h00000000 /* 0x3c28 */;
                3851: data_o = 32'h00000000 /* 0x3c2c */;
                3852: data_o = 32'h00000000 /* 0x3c30 */;
                3853: data_o = 32'h00000000 /* 0x3c34 */;
                3854: data_o = 32'h00000000 /* 0x3c38 */;
                3855: data_o = 32'h00000000 /* 0x3c3c */;
                3856: data_o = 32'h00000000 /* 0x3c40 */;
                3857: data_o = 32'h00000000 /* 0x3c44 */;
                3858: data_o = 32'h00000000 /* 0x3c48 */;
                3859: data_o = 32'h00000000 /* 0x3c4c */;
                3860: data_o = 32'h00000000 /* 0x3c50 */;
                3861: data_o = 32'h00000000 /* 0x3c54 */;
                3862: data_o = 32'h00000000 /* 0x3c58 */;
                3863: data_o = 32'h00000000 /* 0x3c5c */;
                3864: data_o = 32'h00000000 /* 0x3c60 */;
                3865: data_o = 32'h00000000 /* 0x3c64 */;
                3866: data_o = 32'h00000000 /* 0x3c68 */;
                3867: data_o = 32'h00000000 /* 0x3c6c */;
                3868: data_o = 32'h00000000 /* 0x3c70 */;
                3869: data_o = 32'h00000000 /* 0x3c74 */;
                3870: data_o = 32'h00000000 /* 0x3c78 */;
                3871: data_o = 32'h00000000 /* 0x3c7c */;
                3872: data_o = 32'h00000000 /* 0x3c80 */;
                3873: data_o = 32'h00000000 /* 0x3c84 */;
                3874: data_o = 32'h00000000 /* 0x3c88 */;
                3875: data_o = 32'h00000000 /* 0x3c8c */;
                3876: data_o = 32'h00000000 /* 0x3c90 */;
                3877: data_o = 32'h00000000 /* 0x3c94 */;
                3878: data_o = 32'h00000000 /* 0x3c98 */;
                3879: data_o = 32'h00000000 /* 0x3c9c */;
                3880: data_o = 32'h00000000 /* 0x3ca0 */;
                3881: data_o = 32'h00000000 /* 0x3ca4 */;
                3882: data_o = 32'h00000000 /* 0x3ca8 */;
                3883: data_o = 32'h00000000 /* 0x3cac */;
                3884: data_o = 32'h00000000 /* 0x3cb0 */;
                3885: data_o = 32'h00000000 /* 0x3cb4 */;
                3886: data_o = 32'h00000000 /* 0x3cb8 */;
                3887: data_o = 32'h00000000 /* 0x3cbc */;
                3888: data_o = 32'h00000000 /* 0x3cc0 */;
                3889: data_o = 32'h00000000 /* 0x3cc4 */;
                3890: data_o = 32'h00000000 /* 0x3cc8 */;
                3891: data_o = 32'h00000000 /* 0x3ccc */;
                3892: data_o = 32'h00000000 /* 0x3cd0 */;
                3893: data_o = 32'h00000000 /* 0x3cd4 */;
                3894: data_o = 32'h00000000 /* 0x3cd8 */;
                3895: data_o = 32'h00000000 /* 0x3cdc */;
                3896: data_o = 32'h00000000 /* 0x3ce0 */;
                3897: data_o = 32'h00000000 /* 0x3ce4 */;
                3898: data_o = 32'h00000000 /* 0x3ce8 */;
                3899: data_o = 32'h00000000 /* 0x3cec */;
                3900: data_o = 32'h00000000 /* 0x3cf0 */;
                3901: data_o = 32'h00000000 /* 0x3cf4 */;
                3902: data_o = 32'h00000000 /* 0x3cf8 */;
                3903: data_o = 32'h00000000 /* 0x3cfc */;
                3904: data_o = 32'h00000000 /* 0x3d00 */;
                3905: data_o = 32'h00000000 /* 0x3d04 */;
                3906: data_o = 32'h00000000 /* 0x3d08 */;
                3907: data_o = 32'h00000000 /* 0x3d0c */;
                3908: data_o = 32'h00000000 /* 0x3d10 */;
                3909: data_o = 32'h00000000 /* 0x3d14 */;
                3910: data_o = 32'h00000000 /* 0x3d18 */;
                3911: data_o = 32'h00000000 /* 0x3d1c */;
                3912: data_o = 32'h00000000 /* 0x3d20 */;
                3913: data_o = 32'h00000000 /* 0x3d24 */;
                3914: data_o = 32'h00000000 /* 0x3d28 */;
                3915: data_o = 32'h00000000 /* 0x3d2c */;
                3916: data_o = 32'h00000000 /* 0x3d30 */;
                3917: data_o = 32'h00000000 /* 0x3d34 */;
                3918: data_o = 32'h00000000 /* 0x3d38 */;
                3919: data_o = 32'h00000000 /* 0x3d3c */;
                3920: data_o = 32'h00000000 /* 0x3d40 */;
                3921: data_o = 32'h00000000 /* 0x3d44 */;
                3922: data_o = 32'h00000000 /* 0x3d48 */;
                3923: data_o = 32'h00000000 /* 0x3d4c */;
                3924: data_o = 32'h00000000 /* 0x3d50 */;
                3925: data_o = 32'h00000000 /* 0x3d54 */;
                3926: data_o = 32'h00000000 /* 0x3d58 */;
                3927: data_o = 32'h00000000 /* 0x3d5c */;
                3928: data_o = 32'h00000000 /* 0x3d60 */;
                3929: data_o = 32'h00000000 /* 0x3d64 */;
                3930: data_o = 32'h00000000 /* 0x3d68 */;
                3931: data_o = 32'h00000000 /* 0x3d6c */;
                3932: data_o = 32'h00000000 /* 0x3d70 */;
                3933: data_o = 32'h00000000 /* 0x3d74 */;
                3934: data_o = 32'h00000000 /* 0x3d78 */;
                3935: data_o = 32'h00000000 /* 0x3d7c */;
                3936: data_o = 32'h00000000 /* 0x3d80 */;
                3937: data_o = 32'h00000000 /* 0x3d84 */;
                3938: data_o = 32'h00000000 /* 0x3d88 */;
                3939: data_o = 32'h00000000 /* 0x3d8c */;
                3940: data_o = 32'h00000000 /* 0x3d90 */;
                3941: data_o = 32'h00000000 /* 0x3d94 */;
                3942: data_o = 32'h00000000 /* 0x3d98 */;
                3943: data_o = 32'h00000000 /* 0x3d9c */;
                3944: data_o = 32'h00000000 /* 0x3da0 */;
                3945: data_o = 32'h00000000 /* 0x3da4 */;
                3946: data_o = 32'h00000000 /* 0x3da8 */;
                3947: data_o = 32'h00000000 /* 0x3dac */;
                3948: data_o = 32'h00000000 /* 0x3db0 */;
                3949: data_o = 32'h00000000 /* 0x3db4 */;
                3950: data_o = 32'h00000000 /* 0x3db8 */;
                3951: data_o = 32'h00000000 /* 0x3dbc */;
                3952: data_o = 32'h00000000 /* 0x3dc0 */;
                3953: data_o = 32'h00000000 /* 0x3dc4 */;
                3954: data_o = 32'h00000000 /* 0x3dc8 */;
                3955: data_o = 32'h00000000 /* 0x3dcc */;
                3956: data_o = 32'h00000000 /* 0x3dd0 */;
                3957: data_o = 32'h00000000 /* 0x3dd4 */;
                3958: data_o = 32'h00000000 /* 0x3dd8 */;
                3959: data_o = 32'h00000000 /* 0x3ddc */;
                3960: data_o = 32'h00000000 /* 0x3de0 */;
                3961: data_o = 32'h00000000 /* 0x3de4 */;
                3962: data_o = 32'h00000000 /* 0x3de8 */;
                3963: data_o = 32'h00000000 /* 0x3dec */;
                3964: data_o = 32'h00000000 /* 0x3df0 */;
                3965: data_o = 32'h00000000 /* 0x3df4 */;
                3966: data_o = 32'h00000000 /* 0x3df8 */;
                3967: data_o = 32'h00000000 /* 0x3dfc */;
                3968: data_o = 32'h00000000 /* 0x3e00 */;
                3969: data_o = 32'h00000000 /* 0x3e04 */;
                3970: data_o = 32'h00000000 /* 0x3e08 */;
                3971: data_o = 32'h00000000 /* 0x3e0c */;
                3972: data_o = 32'h00000000 /* 0x3e10 */;
                3973: data_o = 32'h00000000 /* 0x3e14 */;
                3974: data_o = 32'h00000000 /* 0x3e18 */;
                3975: data_o = 32'h00000000 /* 0x3e1c */;
                3976: data_o = 32'h00000000 /* 0x3e20 */;
                3977: data_o = 32'h00000000 /* 0x3e24 */;
                3978: data_o = 32'h00000000 /* 0x3e28 */;
                3979: data_o = 32'h00000000 /* 0x3e2c */;
                3980: data_o = 32'h00000000 /* 0x3e30 */;
                3981: data_o = 32'h00000000 /* 0x3e34 */;
                3982: data_o = 32'h00000000 /* 0x3e38 */;
                3983: data_o = 32'h00000000 /* 0x3e3c */;
                3984: data_o = 32'h00000000 /* 0x3e40 */;
                3985: data_o = 32'h00000000 /* 0x3e44 */;
                3986: data_o = 32'h00000000 /* 0x3e48 */;
                3987: data_o = 32'h00000000 /* 0x3e4c */;
                3988: data_o = 32'h00000000 /* 0x3e50 */;
                3989: data_o = 32'h00000000 /* 0x3e54 */;
                3990: data_o = 32'h00000000 /* 0x3e58 */;
                3991: data_o = 32'h00000000 /* 0x3e5c */;
                3992: data_o = 32'h00000000 /* 0x3e60 */;
                3993: data_o = 32'h00000000 /* 0x3e64 */;
                3994: data_o = 32'h00000000 /* 0x3e68 */;
                3995: data_o = 32'h00000000 /* 0x3e6c */;
                3996: data_o = 32'h00000000 /* 0x3e70 */;
                3997: data_o = 32'h00000000 /* 0x3e74 */;
                3998: data_o = 32'h00000000 /* 0x3e78 */;
                3999: data_o = 32'h00000000 /* 0x3e7c */;
                4000: data_o = 32'h00000000 /* 0x3e80 */;
                4001: data_o = 32'h00000000 /* 0x3e84 */;
                4002: data_o = 32'h00000000 /* 0x3e88 */;
                4003: data_o = 32'h00000000 /* 0x3e8c */;
                4004: data_o = 32'h00000000 /* 0x3e90 */;
                4005: data_o = 32'h00000000 /* 0x3e94 */;
                4006: data_o = 32'h00000000 /* 0x3e98 */;
                4007: data_o = 32'h00000000 /* 0x3e9c */;
                4008: data_o = 32'h00000000 /* 0x3ea0 */;
                4009: data_o = 32'h00000000 /* 0x3ea4 */;
                4010: data_o = 32'h00000000 /* 0x3ea8 */;
                4011: data_o = 32'h00000000 /* 0x3eac */;
                4012: data_o = 32'h00000000 /* 0x3eb0 */;
                4013: data_o = 32'h00000000 /* 0x3eb4 */;
                4014: data_o = 32'h00000000 /* 0x3eb8 */;
                4015: data_o = 32'h00000000 /* 0x3ebc */;
                4016: data_o = 32'h00000000 /* 0x3ec0 */;
                4017: data_o = 32'h00000000 /* 0x3ec4 */;
                4018: data_o = 32'h00000000 /* 0x3ec8 */;
                4019: data_o = 32'h00000000 /* 0x3ecc */;
                4020: data_o = 32'h00000000 /* 0x3ed0 */;
                4021: data_o = 32'h00000000 /* 0x3ed4 */;
                4022: data_o = 32'h00000000 /* 0x3ed8 */;
                4023: data_o = 32'h00000000 /* 0x3edc */;
                4024: data_o = 32'h00000000 /* 0x3ee0 */;
                4025: data_o = 32'h00000000 /* 0x3ee4 */;
                4026: data_o = 32'h00000000 /* 0x3ee8 */;
                4027: data_o = 32'h00000000 /* 0x3eec */;
                4028: data_o = 32'h00000000 /* 0x3ef0 */;
                4029: data_o = 32'h00000000 /* 0x3ef4 */;
                4030: data_o = 32'h00000000 /* 0x3ef8 */;
                4031: data_o = 32'h00000000 /* 0x3efc */;
                4032: data_o = 32'h00000000 /* 0x3f00 */;
                4033: data_o = 32'h00000000 /* 0x3f04 */;
                4034: data_o = 32'h00000000 /* 0x3f08 */;
                4035: data_o = 32'h00000000 /* 0x3f0c */;
                4036: data_o = 32'h00000000 /* 0x3f10 */;
                4037: data_o = 32'h00000000 /* 0x3f14 */;
                4038: data_o = 32'h00000000 /* 0x3f18 */;
                4039: data_o = 32'h00000000 /* 0x3f1c */;
                4040: data_o = 32'h00000000 /* 0x3f20 */;
                4041: data_o = 32'h00000000 /* 0x3f24 */;
                4042: data_o = 32'h00000000 /* 0x3f28 */;
                4043: data_o = 32'h00000000 /* 0x3f2c */;
                4044: data_o = 32'h00000000 /* 0x3f30 */;
                4045: data_o = 32'h00000000 /* 0x3f34 */;
                4046: data_o = 32'h00000000 /* 0x3f38 */;
                4047: data_o = 32'h00000000 /* 0x3f3c */;
                4048: data_o = 32'h00000000 /* 0x3f40 */;
                4049: data_o = 32'h00000000 /* 0x3f44 */;
                4050: data_o = 32'h00000000 /* 0x3f48 */;
                4051: data_o = 32'h00000000 /* 0x3f4c */;
                4052: data_o = 32'h00000000 /* 0x3f50 */;
                4053: data_o = 32'h00000000 /* 0x3f54 */;
                4054: data_o = 32'h00000000 /* 0x3f58 */;
                4055: data_o = 32'h00000000 /* 0x3f5c */;
                4056: data_o = 32'h00000000 /* 0x3f60 */;
                4057: data_o = 32'h00000000 /* 0x3f64 */;
                4058: data_o = 32'h00000000 /* 0x3f68 */;
                4059: data_o = 32'h00000000 /* 0x3f6c */;
                4060: data_o = 32'h00000000 /* 0x3f70 */;
                4061: data_o = 32'h00000000 /* 0x3f74 */;
                4062: data_o = 32'h00000000 /* 0x3f78 */;
                4063: data_o = 32'h00000000 /* 0x3f7c */;
                4064: data_o = 32'h00000000 /* 0x3f80 */;
                4065: data_o = 32'h00000000 /* 0x3f84 */;
                4066: data_o = 32'h00000000 /* 0x3f88 */;
                4067: data_o = 32'h00000000 /* 0x3f8c */;
                4068: data_o = 32'h00000000 /* 0x3f90 */;
                4069: data_o = 32'h00000000 /* 0x3f94 */;
                4070: data_o = 32'h00000000 /* 0x3f98 */;
                4071: data_o = 32'h00000000 /* 0x3f9c */;
                4072: data_o = 32'h00000000 /* 0x3fa0 */;
                4073: data_o = 32'h00000000 /* 0x3fa4 */;
                4074: data_o = 32'h00000000 /* 0x3fa8 */;
                4075: data_o = 32'h00000000 /* 0x3fac */;
                4076: data_o = 32'h00000000 /* 0x3fb0 */;
                4077: data_o = 32'h00000000 /* 0x3fb4 */;
                4078: data_o = 32'h00000000 /* 0x3fb8 */;
                4079: data_o = 32'h00000000 /* 0x3fbc */;
                4080: data_o = 32'h00000000 /* 0x3fc0 */;
                4081: data_o = 32'h00000000 /* 0x3fc4 */;
                4082: data_o = 32'h00000000 /* 0x3fc8 */;
                4083: data_o = 32'h00000000 /* 0x3fcc */;
                4084: data_o = 32'h00000000 /* 0x3fd0 */;
                4085: data_o = 32'h00000000 /* 0x3fd4 */;
                4086: data_o = 32'h00000000 /* 0x3fd8 */;
                4087: data_o = 32'h00000000 /* 0x3fdc */;
                4088: data_o = 32'h00000000 /* 0x3fe0 */;
                4089: data_o = 32'h00000000 /* 0x3fe4 */;
                4090: data_o = 32'h00000000 /* 0x3fe8 */;
                4091: data_o = 32'h00000000 /* 0x3fec */;
                4092: data_o = 32'h00000000 /* 0x3ff0 */;
                4093: data_o = 32'h00000000 /* 0x3ff4 */;
                4094: data_o = 32'h00000000 /* 0x3ff8 */;
                4095: data_o = 32'h00000000 /* 0x3ffc */;
                4096: data_o = 32'h00000000 /* 0x4000 */;
                4097: data_o = 32'h00000000 /* 0x4004 */;
                4098: data_o = 32'h00000000 /* 0x4008 */;
                4099: data_o = 32'h00000000 /* 0x400c */;
                4100: data_o = 32'h00000000 /* 0x4010 */;
                4101: data_o = 32'h00000000 /* 0x4014 */;
                4102: data_o = 32'h00000000 /* 0x4018 */;
                4103: data_o = 32'h00000000 /* 0x401c */;
                4104: data_o = 32'h00000000 /* 0x4020 */;
                4105: data_o = 32'h00000000 /* 0x4024 */;
                4106: data_o = 32'h00000000 /* 0x4028 */;
                4107: data_o = 32'h00000000 /* 0x402c */;
                4108: data_o = 32'h00000000 /* 0x4030 */;
                4109: data_o = 32'h00000000 /* 0x4034 */;
                4110: data_o = 32'h00000000 /* 0x4038 */;
                4111: data_o = 32'h00000000 /* 0x403c */;
                4112: data_o = 32'h00000000 /* 0x4040 */;
                4113: data_o = 32'h00000000 /* 0x4044 */;
                4114: data_o = 32'h00000000 /* 0x4048 */;
                4115: data_o = 32'h00000000 /* 0x404c */;
                4116: data_o = 32'h00000000 /* 0x4050 */;
                4117: data_o = 32'h00000000 /* 0x4054 */;
                4118: data_o = 32'h00000000 /* 0x4058 */;
                4119: data_o = 32'h00000000 /* 0x405c */;
                4120: data_o = 32'h00000000 /* 0x4060 */;
                4121: data_o = 32'h00000000 /* 0x4064 */;
                4122: data_o = 32'h00000000 /* 0x4068 */;
                4123: data_o = 32'h00000000 /* 0x406c */;
                4124: data_o = 32'h00000000 /* 0x4070 */;
                4125: data_o = 32'h00000000 /* 0x4074 */;
                4126: data_o = 32'h00000000 /* 0x4078 */;
                4127: data_o = 32'h00000000 /* 0x407c */;
                4128: data_o = 32'h00000000 /* 0x4080 */;
                4129: data_o = 32'h00000000 /* 0x4084 */;
                4130: data_o = 32'h00000000 /* 0x4088 */;
                4131: data_o = 32'h00000000 /* 0x408c */;
                4132: data_o = 32'h00000000 /* 0x4090 */;
                4133: data_o = 32'h00000000 /* 0x4094 */;
                4134: data_o = 32'h00000000 /* 0x4098 */;
                4135: data_o = 32'h00000000 /* 0x409c */;
                4136: data_o = 32'h00000000 /* 0x40a0 */;
                4137: data_o = 32'h00000000 /* 0x40a4 */;
                4138: data_o = 32'h00000000 /* 0x40a8 */;
                4139: data_o = 32'h00000000 /* 0x40ac */;
                4140: data_o = 32'h00000000 /* 0x40b0 */;
                4141: data_o = 32'h00000000 /* 0x40b4 */;
                4142: data_o = 32'h00000000 /* 0x40b8 */;
                4143: data_o = 32'h00000000 /* 0x40bc */;
                4144: data_o = 32'h00000000 /* 0x40c0 */;
                4145: data_o = 32'h00000000 /* 0x40c4 */;
                4146: data_o = 32'h00000000 /* 0x40c8 */;
                4147: data_o = 32'h00000000 /* 0x40cc */;
                4148: data_o = 32'h00000000 /* 0x40d0 */;
                4149: data_o = 32'h00000000 /* 0x40d4 */;
                4150: data_o = 32'h00000000 /* 0x40d8 */;
                4151: data_o = 32'h00000000 /* 0x40dc */;
                4152: data_o = 32'h00000000 /* 0x40e0 */;
                4153: data_o = 32'h00000000 /* 0x40e4 */;
                4154: data_o = 32'h00000000 /* 0x40e8 */;
                4155: data_o = 32'h00000000 /* 0x40ec */;
                4156: data_o = 32'h00000000 /* 0x40f0 */;
                4157: data_o = 32'h00000000 /* 0x40f4 */;
                4158: data_o = 32'h00000000 /* 0x40f8 */;
                4159: data_o = 32'h00000000 /* 0x40fc */;
                4160: data_o = 32'h00000000 /* 0x4100 */;
                4161: data_o = 32'h00000000 /* 0x4104 */;
                4162: data_o = 32'h00000000 /* 0x4108 */;
                4163: data_o = 32'h00000000 /* 0x410c */;
                4164: data_o = 32'h00000000 /* 0x4110 */;
                4165: data_o = 32'h00000000 /* 0x4114 */;
                4166: data_o = 32'h00000000 /* 0x4118 */;
                4167: data_o = 32'h00000000 /* 0x411c */;
                4168: data_o = 32'h00000000 /* 0x4120 */;
                4169: data_o = 32'h00000000 /* 0x4124 */;
                4170: data_o = 32'h00000000 /* 0x4128 */;
                4171: data_o = 32'h00000000 /* 0x412c */;
                4172: data_o = 32'h00000000 /* 0x4130 */;
                4173: data_o = 32'h00000000 /* 0x4134 */;
                4174: data_o = 32'h00000000 /* 0x4138 */;
                4175: data_o = 32'h00000000 /* 0x413c */;
                4176: data_o = 32'h00000000 /* 0x4140 */;
                4177: data_o = 32'h00000000 /* 0x4144 */;
                4178: data_o = 32'h00000000 /* 0x4148 */;
                4179: data_o = 32'h00000000 /* 0x414c */;
                4180: data_o = 32'h00000000 /* 0x4150 */;
                4181: data_o = 32'h00000000 /* 0x4154 */;
                4182: data_o = 32'h00000000 /* 0x4158 */;
                4183: data_o = 32'h00000000 /* 0x415c */;
                4184: data_o = 32'h00000000 /* 0x4160 */;
                4185: data_o = 32'h00000000 /* 0x4164 */;
                4186: data_o = 32'h00000000 /* 0x4168 */;
                4187: data_o = 32'h00000000 /* 0x416c */;
                4188: data_o = 32'h00000000 /* 0x4170 */;
                4189: data_o = 32'h00000000 /* 0x4174 */;
                4190: data_o = 32'h00000000 /* 0x4178 */;
                4191: data_o = 32'h00000000 /* 0x417c */;
                4192: data_o = 32'h00000000 /* 0x4180 */;
                4193: data_o = 32'h00000000 /* 0x4184 */;
                4194: data_o = 32'h00000000 /* 0x4188 */;
                4195: data_o = 32'h00000000 /* 0x418c */;
                4196: data_o = 32'h00000000 /* 0x4190 */;
                4197: data_o = 32'h00000000 /* 0x4194 */;
                4198: data_o = 32'h00000000 /* 0x4198 */;
                4199: data_o = 32'h00000000 /* 0x419c */;
                4200: data_o = 32'h00000000 /* 0x41a0 */;
                4201: data_o = 32'h00000000 /* 0x41a4 */;
                4202: data_o = 32'h00000000 /* 0x41a8 */;
                4203: data_o = 32'h00000000 /* 0x41ac */;
                4204: data_o = 32'h00000000 /* 0x41b0 */;
                4205: data_o = 32'h00000000 /* 0x41b4 */;
                4206: data_o = 32'h00000000 /* 0x41b8 */;
                4207: data_o = 32'h00000000 /* 0x41bc */;
                4208: data_o = 32'h00000000 /* 0x41c0 */;
                4209: data_o = 32'h00000000 /* 0x41c4 */;
                4210: data_o = 32'h00000000 /* 0x41c8 */;
                4211: data_o = 32'h00000000 /* 0x41cc */;
                4212: data_o = 32'h00000000 /* 0x41d0 */;
                4213: data_o = 32'h00000000 /* 0x41d4 */;
                4214: data_o = 32'h00000000 /* 0x41d8 */;
                4215: data_o = 32'h00000000 /* 0x41dc */;
                4216: data_o = 32'h00000000 /* 0x41e0 */;
                4217: data_o = 32'h00000000 /* 0x41e4 */;
                4218: data_o = 32'h00000000 /* 0x41e8 */;
                4219: data_o = 32'h00000000 /* 0x41ec */;
                4220: data_o = 32'h00000000 /* 0x41f0 */;
                4221: data_o = 32'h00000000 /* 0x41f4 */;
                4222: data_o = 32'h00000000 /* 0x41f8 */;
                4223: data_o = 32'h00000000 /* 0x41fc */;
                4224: data_o = 32'h00000000 /* 0x4200 */;
                4225: data_o = 32'h00000000 /* 0x4204 */;
                4226: data_o = 32'h00000000 /* 0x4208 */;
                4227: data_o = 32'h00000000 /* 0x420c */;
                4228: data_o = 32'h00000000 /* 0x4210 */;
                4229: data_o = 32'h00000000 /* 0x4214 */;
                4230: data_o = 32'h00000000 /* 0x4218 */;
                4231: data_o = 32'h00000000 /* 0x421c */;
                4232: data_o = 32'h00000000 /* 0x4220 */;
                4233: data_o = 32'h00000000 /* 0x4224 */;
                4234: data_o = 32'h00000000 /* 0x4228 */;
                4235: data_o = 32'h00000000 /* 0x422c */;
                4236: data_o = 32'h00000000 /* 0x4230 */;
                4237: data_o = 32'h00000000 /* 0x4234 */;
                4238: data_o = 32'h00000000 /* 0x4238 */;
                4239: data_o = 32'h00000000 /* 0x423c */;
                4240: data_o = 32'h00000000 /* 0x4240 */;
                4241: data_o = 32'h00000000 /* 0x4244 */;
                4242: data_o = 32'h00000000 /* 0x4248 */;
                4243: data_o = 32'h00000000 /* 0x424c */;
                4244: data_o = 32'h00000000 /* 0x4250 */;
                4245: data_o = 32'h00000000 /* 0x4254 */;
                4246: data_o = 32'h00000000 /* 0x4258 */;
                4247: data_o = 32'h00000000 /* 0x425c */;
                4248: data_o = 32'h00000000 /* 0x4260 */;
                4249: data_o = 32'h00000000 /* 0x4264 */;
                4250: data_o = 32'h00000000 /* 0x4268 */;
                4251: data_o = 32'h00000000 /* 0x426c */;
                4252: data_o = 32'h00000000 /* 0x4270 */;
                4253: data_o = 32'h00000000 /* 0x4274 */;
                4254: data_o = 32'h00000000 /* 0x4278 */;
                4255: data_o = 32'h00000000 /* 0x427c */;
                4256: data_o = 32'h00000000 /* 0x4280 */;
                4257: data_o = 32'h00000000 /* 0x4284 */;
                4258: data_o = 32'h00000000 /* 0x4288 */;
                4259: data_o = 32'h00000000 /* 0x428c */;
                4260: data_o = 32'h00000000 /* 0x4290 */;
                4261: data_o = 32'h00000000 /* 0x4294 */;
                4262: data_o = 32'h00000000 /* 0x4298 */;
                4263: data_o = 32'h00000000 /* 0x429c */;
                4264: data_o = 32'h00000000 /* 0x42a0 */;
                4265: data_o = 32'h00000000 /* 0x42a4 */;
                4266: data_o = 32'h00000000 /* 0x42a8 */;
                4267: data_o = 32'h00000000 /* 0x42ac */;
                4268: data_o = 32'h00000000 /* 0x42b0 */;
                4269: data_o = 32'h00000000 /* 0x42b4 */;
                4270: data_o = 32'h00000000 /* 0x42b8 */;
                4271: data_o = 32'h00000000 /* 0x42bc */;
                4272: data_o = 32'h00000000 /* 0x42c0 */;
                4273: data_o = 32'h00000000 /* 0x42c4 */;
                4274: data_o = 32'h00000000 /* 0x42c8 */;
                4275: data_o = 32'h00000000 /* 0x42cc */;
                4276: data_o = 32'h00000000 /* 0x42d0 */;
                4277: data_o = 32'h00000000 /* 0x42d4 */;
                4278: data_o = 32'h00000000 /* 0x42d8 */;
                4279: data_o = 32'h00000000 /* 0x42dc */;
                4280: data_o = 32'h00000000 /* 0x42e0 */;
                4281: data_o = 32'h00000000 /* 0x42e4 */;
                4282: data_o = 32'h00000000 /* 0x42e8 */;
                4283: data_o = 32'h00000000 /* 0x42ec */;
                4284: data_o = 32'h00000000 /* 0x42f0 */;
                4285: data_o = 32'h00000000 /* 0x42f4 */;
                4286: data_o = 32'h00000000 /* 0x42f8 */;
                4287: data_o = 32'h00000000 /* 0x42fc */;
                4288: data_o = 32'h00000000 /* 0x4300 */;
                4289: data_o = 32'h00000000 /* 0x4304 */;
                4290: data_o = 32'h00000000 /* 0x4308 */;
                4291: data_o = 32'h00000000 /* 0x430c */;
                4292: data_o = 32'h00000000 /* 0x4310 */;
                4293: data_o = 32'h00000000 /* 0x4314 */;
                4294: data_o = 32'h00000000 /* 0x4318 */;
                4295: data_o = 32'h00000000 /* 0x431c */;
                4296: data_o = 32'h00000000 /* 0x4320 */;
                4297: data_o = 32'h00000000 /* 0x4324 */;
                4298: data_o = 32'h00000000 /* 0x4328 */;
                4299: data_o = 32'h00000000 /* 0x432c */;
                4300: data_o = 32'h00000000 /* 0x4330 */;
                4301: data_o = 32'h00000000 /* 0x4334 */;
                4302: data_o = 32'h00000000 /* 0x4338 */;
                4303: data_o = 32'h00000000 /* 0x433c */;
                4304: data_o = 32'h00000000 /* 0x4340 */;
                4305: data_o = 32'h00000000 /* 0x4344 */;
                4306: data_o = 32'h00000000 /* 0x4348 */;
                4307: data_o = 32'h00000000 /* 0x434c */;
                4308: data_o = 32'h00000000 /* 0x4350 */;
                4309: data_o = 32'h00000000 /* 0x4354 */;
                4310: data_o = 32'h00000000 /* 0x4358 */;
                4311: data_o = 32'h00000000 /* 0x435c */;
                4312: data_o = 32'h00000000 /* 0x4360 */;
                4313: data_o = 32'h00000000 /* 0x4364 */;
                4314: data_o = 32'h00000000 /* 0x4368 */;
                4315: data_o = 32'h00000000 /* 0x436c */;
                4316: data_o = 32'h00000000 /* 0x4370 */;
                4317: data_o = 32'h00000000 /* 0x4374 */;
                4318: data_o = 32'h00000000 /* 0x4378 */;
                4319: data_o = 32'h00000000 /* 0x437c */;
                4320: data_o = 32'h00000000 /* 0x4380 */;
                4321: data_o = 32'h00000000 /* 0x4384 */;
                4322: data_o = 32'h00000000 /* 0x4388 */;
                4323: data_o = 32'h00000000 /* 0x438c */;
                4324: data_o = 32'h00000000 /* 0x4390 */;
                4325: data_o = 32'h00000000 /* 0x4394 */;
                4326: data_o = 32'h00000000 /* 0x4398 */;
                4327: data_o = 32'h00000000 /* 0x439c */;
                4328: data_o = 32'h00000000 /* 0x43a0 */;
                4329: data_o = 32'h00000000 /* 0x43a4 */;
                4330: data_o = 32'h00000000 /* 0x43a8 */;
                4331: data_o = 32'h00000000 /* 0x43ac */;
                4332: data_o = 32'h00000000 /* 0x43b0 */;
                4333: data_o = 32'h00000000 /* 0x43b4 */;
                4334: data_o = 32'h00000000 /* 0x43b8 */;
                4335: data_o = 32'h00000000 /* 0x43bc */;
                4336: data_o = 32'h00000000 /* 0x43c0 */;
                4337: data_o = 32'h00000000 /* 0x43c4 */;
                4338: data_o = 32'h00000000 /* 0x43c8 */;
                4339: data_o = 32'h00000000 /* 0x43cc */;
                4340: data_o = 32'h00000000 /* 0x43d0 */;
                4341: data_o = 32'h00000000 /* 0x43d4 */;
                4342: data_o = 32'h00000000 /* 0x43d8 */;
                4343: data_o = 32'h00000000 /* 0x43dc */;
                4344: data_o = 32'h00000000 /* 0x43e0 */;
                4345: data_o = 32'h00000000 /* 0x43e4 */;
                4346: data_o = 32'h00000000 /* 0x43e8 */;
                4347: data_o = 32'h00000000 /* 0x43ec */;
                4348: data_o = 32'h00000000 /* 0x43f0 */;
                4349: data_o = 32'h00000000 /* 0x43f4 */;
                4350: data_o = 32'h00000000 /* 0x43f8 */;
                4351: data_o = 32'h00000000 /* 0x43fc */;
                4352: data_o = 32'h00000000 /* 0x4400 */;
                4353: data_o = 32'h00000000 /* 0x4404 */;
                4354: data_o = 32'h00000000 /* 0x4408 */;
                4355: data_o = 32'h00000000 /* 0x440c */;
                4356: data_o = 32'h00000000 /* 0x4410 */;
                4357: data_o = 32'h00000000 /* 0x4414 */;
                4358: data_o = 32'h00000000 /* 0x4418 */;
                4359: data_o = 32'h00000000 /* 0x441c */;
                4360: data_o = 32'h00000000 /* 0x4420 */;
                4361: data_o = 32'h00000000 /* 0x4424 */;
                4362: data_o = 32'h00000000 /* 0x4428 */;
                4363: data_o = 32'h00000000 /* 0x442c */;
                4364: data_o = 32'h00000000 /* 0x4430 */;
                4365: data_o = 32'h00000000 /* 0x4434 */;
                4366: data_o = 32'h00000000 /* 0x4438 */;
                4367: data_o = 32'h00000000 /* 0x443c */;
                4368: data_o = 32'h00000000 /* 0x4440 */;
                4369: data_o = 32'h00000000 /* 0x4444 */;
                4370: data_o = 32'h00000000 /* 0x4448 */;
                4371: data_o = 32'h00000000 /* 0x444c */;
                4372: data_o = 32'h00000000 /* 0x4450 */;
                4373: data_o = 32'h00000000 /* 0x4454 */;
                4374: data_o = 32'h00000000 /* 0x4458 */;
                4375: data_o = 32'h00000000 /* 0x445c */;
                4376: data_o = 32'h00000000 /* 0x4460 */;
                4377: data_o = 32'h00000000 /* 0x4464 */;
                4378: data_o = 32'h00000000 /* 0x4468 */;
                4379: data_o = 32'h00000000 /* 0x446c */;
                4380: data_o = 32'h00000000 /* 0x4470 */;
                4381: data_o = 32'h00000000 /* 0x4474 */;
                4382: data_o = 32'h00000000 /* 0x4478 */;
                4383: data_o = 32'h00000000 /* 0x447c */;
                4384: data_o = 32'h00000000 /* 0x4480 */;
                4385: data_o = 32'h00000000 /* 0x4484 */;
                4386: data_o = 32'h00000000 /* 0x4488 */;
                4387: data_o = 32'h00000000 /* 0x448c */;
                4388: data_o = 32'h00000000 /* 0x4490 */;
                4389: data_o = 32'h00000000 /* 0x4494 */;
                4390: data_o = 32'h00000000 /* 0x4498 */;
                4391: data_o = 32'h00000000 /* 0x449c */;
                4392: data_o = 32'h00000000 /* 0x44a0 */;
                4393: data_o = 32'h00000000 /* 0x44a4 */;
                4394: data_o = 32'h00000000 /* 0x44a8 */;
                4395: data_o = 32'h00000000 /* 0x44ac */;
                4396: data_o = 32'h00000000 /* 0x44b0 */;
                4397: data_o = 32'h00000000 /* 0x44b4 */;
                4398: data_o = 32'h00000000 /* 0x44b8 */;
                4399: data_o = 32'h00000000 /* 0x44bc */;
                4400: data_o = 32'h00000000 /* 0x44c0 */;
                4401: data_o = 32'h00000000 /* 0x44c4 */;
                4402: data_o = 32'h00000000 /* 0x44c8 */;
                4403: data_o = 32'h00000000 /* 0x44cc */;
                4404: data_o = 32'h00000000 /* 0x44d0 */;
                4405: data_o = 32'h00000000 /* 0x44d4 */;
                4406: data_o = 32'h00000000 /* 0x44d8 */;
                4407: data_o = 32'h00000000 /* 0x44dc */;
                4408: data_o = 32'h00000000 /* 0x44e0 */;
                4409: data_o = 32'h00000000 /* 0x44e4 */;
                4410: data_o = 32'h00000000 /* 0x44e8 */;
                4411: data_o = 32'h00000000 /* 0x44ec */;
                4412: data_o = 32'h00000000 /* 0x44f0 */;
                4413: data_o = 32'h00000000 /* 0x44f4 */;
                4414: data_o = 32'h00000000 /* 0x44f8 */;
                4415: data_o = 32'h00000000 /* 0x44fc */;
                4416: data_o = 32'h00000000 /* 0x4500 */;
                4417: data_o = 32'h00000000 /* 0x4504 */;
                4418: data_o = 32'h00000000 /* 0x4508 */;
                4419: data_o = 32'h00000000 /* 0x450c */;
                4420: data_o = 32'h00000000 /* 0x4510 */;
                4421: data_o = 32'h00000000 /* 0x4514 */;
                4422: data_o = 32'h00000000 /* 0x4518 */;
                4423: data_o = 32'h00000000 /* 0x451c */;
                4424: data_o = 32'h00000000 /* 0x4520 */;
                4425: data_o = 32'h00000000 /* 0x4524 */;
                4426: data_o = 32'h00000000 /* 0x4528 */;
                4427: data_o = 32'h00000000 /* 0x452c */;
                4428: data_o = 32'h00000000 /* 0x4530 */;
                4429: data_o = 32'h00000000 /* 0x4534 */;
                4430: data_o = 32'h00000000 /* 0x4538 */;
                4431: data_o = 32'h00000000 /* 0x453c */;
                4432: data_o = 32'h00000000 /* 0x4540 */;
                4433: data_o = 32'h00000000 /* 0x4544 */;
                4434: data_o = 32'h00000000 /* 0x4548 */;
                4435: data_o = 32'h00000000 /* 0x454c */;
                4436: data_o = 32'h00000000 /* 0x4550 */;
                4437: data_o = 32'h00000000 /* 0x4554 */;
                4438: data_o = 32'h00000000 /* 0x4558 */;
                4439: data_o = 32'h00000000 /* 0x455c */;
                4440: data_o = 32'h00000000 /* 0x4560 */;
                4441: data_o = 32'h00000000 /* 0x4564 */;
                4442: data_o = 32'h00000000 /* 0x4568 */;
                4443: data_o = 32'h00000000 /* 0x456c */;
                4444: data_o = 32'h00000000 /* 0x4570 */;
                4445: data_o = 32'h00000000 /* 0x4574 */;
                4446: data_o = 32'h00000000 /* 0x4578 */;
                4447: data_o = 32'h00000000 /* 0x457c */;
                4448: data_o = 32'h00000000 /* 0x4580 */;
                4449: data_o = 32'h00000000 /* 0x4584 */;
                4450: data_o = 32'h00000000 /* 0x4588 */;
                4451: data_o = 32'h00000000 /* 0x458c */;
                4452: data_o = 32'h00000000 /* 0x4590 */;
                4453: data_o = 32'h00000000 /* 0x4594 */;
                4454: data_o = 32'h00000000 /* 0x4598 */;
                4455: data_o = 32'h00000000 /* 0x459c */;
                4456: data_o = 32'h00000000 /* 0x45a0 */;
                4457: data_o = 32'h00000000 /* 0x45a4 */;
                4458: data_o = 32'h00000000 /* 0x45a8 */;
                4459: data_o = 32'h00000000 /* 0x45ac */;
                4460: data_o = 32'h00000000 /* 0x45b0 */;
                4461: data_o = 32'h00000000 /* 0x45b4 */;
                4462: data_o = 32'h00000000 /* 0x45b8 */;
                4463: data_o = 32'h00000000 /* 0x45bc */;
                4464: data_o = 32'h00000000 /* 0x45c0 */;
                4465: data_o = 32'h00000000 /* 0x45c4 */;
                4466: data_o = 32'h00000000 /* 0x45c8 */;
                4467: data_o = 32'h00000000 /* 0x45cc */;
                4468: data_o = 32'h00000000 /* 0x45d0 */;
                4469: data_o = 32'h00000000 /* 0x45d4 */;
                4470: data_o = 32'h00000000 /* 0x45d8 */;
                4471: data_o = 32'h00000000 /* 0x45dc */;
                4472: data_o = 32'h00000000 /* 0x45e0 */;
                4473: data_o = 32'h00000000 /* 0x45e4 */;
                4474: data_o = 32'h00000000 /* 0x45e8 */;
                4475: data_o = 32'h00000000 /* 0x45ec */;
                4476: data_o = 32'h00000000 /* 0x45f0 */;
                4477: data_o = 32'h00000000 /* 0x45f4 */;
                4478: data_o = 32'h00000000 /* 0x45f8 */;
                4479: data_o = 32'h00000000 /* 0x45fc */;
                4480: data_o = 32'h00000000 /* 0x4600 */;
                4481: data_o = 32'h00000000 /* 0x4604 */;
                4482: data_o = 32'h00000000 /* 0x4608 */;
                4483: data_o = 32'h00000000 /* 0x460c */;
                4484: data_o = 32'h00000000 /* 0x4610 */;
                4485: data_o = 32'h00000000 /* 0x4614 */;
                4486: data_o = 32'h00000000 /* 0x4618 */;
                4487: data_o = 32'h00000000 /* 0x461c */;
                4488: data_o = 32'h00000000 /* 0x4620 */;
                4489: data_o = 32'h00000000 /* 0x4624 */;
                4490: data_o = 32'h00000000 /* 0x4628 */;
                4491: data_o = 32'h00000000 /* 0x462c */;
                4492: data_o = 32'h00000000 /* 0x4630 */;
                4493: data_o = 32'h00000000 /* 0x4634 */;
                4494: data_o = 32'h00000000 /* 0x4638 */;
                4495: data_o = 32'h00000000 /* 0x463c */;
                4496: data_o = 32'h00000000 /* 0x4640 */;
                4497: data_o = 32'h00000000 /* 0x4644 */;
                4498: data_o = 32'h00000000 /* 0x4648 */;
                4499: data_o = 32'h00000000 /* 0x464c */;
                4500: data_o = 32'h00000000 /* 0x4650 */;
                4501: data_o = 32'h00000000 /* 0x4654 */;
                4502: data_o = 32'h00000000 /* 0x4658 */;
                4503: data_o = 32'h00000000 /* 0x465c */;
                4504: data_o = 32'h00000000 /* 0x4660 */;
                4505: data_o = 32'h00000000 /* 0x4664 */;
                4506: data_o = 32'h00000000 /* 0x4668 */;
                4507: data_o = 32'h00000000 /* 0x466c */;
                4508: data_o = 32'h00000000 /* 0x4670 */;
                4509: data_o = 32'h00000000 /* 0x4674 */;
                4510: data_o = 32'h00000000 /* 0x4678 */;
                4511: data_o = 32'h00000000 /* 0x467c */;
                4512: data_o = 32'h00000000 /* 0x4680 */;
                4513: data_o = 32'h00000000 /* 0x4684 */;
                4514: data_o = 32'h00000000 /* 0x4688 */;
                4515: data_o = 32'h00000000 /* 0x468c */;
                4516: data_o = 32'h00000000 /* 0x4690 */;
                4517: data_o = 32'h00000000 /* 0x4694 */;
                4518: data_o = 32'h00000000 /* 0x4698 */;
                4519: data_o = 32'h00000000 /* 0x469c */;
                4520: data_o = 32'h00000000 /* 0x46a0 */;
                4521: data_o = 32'h00000000 /* 0x46a4 */;
                4522: data_o = 32'h00000000 /* 0x46a8 */;
                4523: data_o = 32'h00000000 /* 0x46ac */;
                4524: data_o = 32'h00000000 /* 0x46b0 */;
                4525: data_o = 32'h00000000 /* 0x46b4 */;
                4526: data_o = 32'h00000000 /* 0x46b8 */;
                4527: data_o = 32'h00000000 /* 0x46bc */;
                4528: data_o = 32'h00000000 /* 0x46c0 */;
                4529: data_o = 32'h00000000 /* 0x46c4 */;
                4530: data_o = 32'h00000000 /* 0x46c8 */;
                4531: data_o = 32'h00000000 /* 0x46cc */;
                4532: data_o = 32'h00000000 /* 0x46d0 */;
                4533: data_o = 32'h00000000 /* 0x46d4 */;
                4534: data_o = 32'h00000000 /* 0x46d8 */;
                4535: data_o = 32'h00000000 /* 0x46dc */;
                4536: data_o = 32'h00000000 /* 0x46e0 */;
                4537: data_o = 32'h00000000 /* 0x46e4 */;
                4538: data_o = 32'h00000000 /* 0x46e8 */;
                4539: data_o = 32'h00000000 /* 0x46ec */;
                4540: data_o = 32'h00000000 /* 0x46f0 */;
                4541: data_o = 32'h00000000 /* 0x46f4 */;
                4542: data_o = 32'h00000000 /* 0x46f8 */;
                4543: data_o = 32'h00000000 /* 0x46fc */;
                4544: data_o = 32'h00000000 /* 0x4700 */;
                4545: data_o = 32'h00000000 /* 0x4704 */;
                4546: data_o = 32'h00000000 /* 0x4708 */;
                4547: data_o = 32'h00000000 /* 0x470c */;
                4548: data_o = 32'h00000000 /* 0x4710 */;
                4549: data_o = 32'h00000000 /* 0x4714 */;
                4550: data_o = 32'h00000000 /* 0x4718 */;
                4551: data_o = 32'h00000000 /* 0x471c */;
                4552: data_o = 32'h00000000 /* 0x4720 */;
                4553: data_o = 32'h00000000 /* 0x4724 */;
                4554: data_o = 32'h00000000 /* 0x4728 */;
                4555: data_o = 32'h00000000 /* 0x472c */;
                4556: data_o = 32'h00000000 /* 0x4730 */;
                4557: data_o = 32'h00000000 /* 0x4734 */;
                4558: data_o = 32'h00000000 /* 0x4738 */;
                4559: data_o = 32'h00000000 /* 0x473c */;
                4560: data_o = 32'h00000000 /* 0x4740 */;
                4561: data_o = 32'h00000000 /* 0x4744 */;
                4562: data_o = 32'h00000000 /* 0x4748 */;
                4563: data_o = 32'h00000000 /* 0x474c */;
                4564: data_o = 32'h00000000 /* 0x4750 */;
                4565: data_o = 32'h00000000 /* 0x4754 */;
                4566: data_o = 32'h00000000 /* 0x4758 */;
                4567: data_o = 32'h00000000 /* 0x475c */;
                4568: data_o = 32'h00000000 /* 0x4760 */;
                4569: data_o = 32'h00000000 /* 0x4764 */;
                4570: data_o = 32'h00000000 /* 0x4768 */;
                4571: data_o = 32'h00000000 /* 0x476c */;
                4572: data_o = 32'h00000000 /* 0x4770 */;
                4573: data_o = 32'h00000000 /* 0x4774 */;
                4574: data_o = 32'h00000000 /* 0x4778 */;
                4575: data_o = 32'h00000000 /* 0x477c */;
                4576: data_o = 32'h00000000 /* 0x4780 */;
                4577: data_o = 32'h00000000 /* 0x4784 */;
                4578: data_o = 32'h00000000 /* 0x4788 */;
                4579: data_o = 32'h00000000 /* 0x478c */;
                4580: data_o = 32'h00000000 /* 0x4790 */;
                4581: data_o = 32'h00000000 /* 0x4794 */;
                4582: data_o = 32'h00000000 /* 0x4798 */;
                4583: data_o = 32'h00000000 /* 0x479c */;
                4584: data_o = 32'h00000000 /* 0x47a0 */;
                4585: data_o = 32'h00000000 /* 0x47a4 */;
                4586: data_o = 32'h00000000 /* 0x47a8 */;
                4587: data_o = 32'h00000000 /* 0x47ac */;
                4588: data_o = 32'h00000000 /* 0x47b0 */;
                4589: data_o = 32'h00000000 /* 0x47b4 */;
                4590: data_o = 32'h00000000 /* 0x47b8 */;
                4591: data_o = 32'h00000000 /* 0x47bc */;
                4592: data_o = 32'h00000000 /* 0x47c0 */;
                4593: data_o = 32'h00000000 /* 0x47c4 */;
                4594: data_o = 32'h00000000 /* 0x47c8 */;
                4595: data_o = 32'h00000000 /* 0x47cc */;
                4596: data_o = 32'h00000000 /* 0x47d0 */;
                4597: data_o = 32'h00000000 /* 0x47d4 */;
                4598: data_o = 32'h00000000 /* 0x47d8 */;
                4599: data_o = 32'h00000000 /* 0x47dc */;
                4600: data_o = 32'h00000000 /* 0x47e0 */;
                4601: data_o = 32'h00000000 /* 0x47e4 */;
                4602: data_o = 32'h00000000 /* 0x47e8 */;
                4603: data_o = 32'h00000000 /* 0x47ec */;
                4604: data_o = 32'h00000000 /* 0x47f0 */;
                4605: data_o = 32'h00000000 /* 0x47f4 */;
                4606: data_o = 32'h00000000 /* 0x47f8 */;
                4607: data_o = 32'h00000000 /* 0x47fc */;
                4608: data_o = 32'h00000000 /* 0x4800 */;
                4609: data_o = 32'h00000000 /* 0x4804 */;
                4610: data_o = 32'h00000000 /* 0x4808 */;
                4611: data_o = 32'h00000000 /* 0x480c */;
                4612: data_o = 32'h00000000 /* 0x4810 */;
                4613: data_o = 32'h00000000 /* 0x4814 */;
                4614: data_o = 32'h00000000 /* 0x4818 */;
                4615: data_o = 32'h00000000 /* 0x481c */;
                4616: data_o = 32'h00000000 /* 0x4820 */;
                4617: data_o = 32'h00000000 /* 0x4824 */;
                4618: data_o = 32'h00000000 /* 0x4828 */;
                4619: data_o = 32'h00000000 /* 0x482c */;
                4620: data_o = 32'h00000000 /* 0x4830 */;
                4621: data_o = 32'h00000000 /* 0x4834 */;
                4622: data_o = 32'h00000000 /* 0x4838 */;
                4623: data_o = 32'h00000000 /* 0x483c */;
                4624: data_o = 32'h00000000 /* 0x4840 */;
                4625: data_o = 32'h00000000 /* 0x4844 */;
                4626: data_o = 32'h00000000 /* 0x4848 */;
                4627: data_o = 32'h00000000 /* 0x484c */;
                4628: data_o = 32'h00000000 /* 0x4850 */;
                4629: data_o = 32'h00000000 /* 0x4854 */;
                4630: data_o = 32'h00000000 /* 0x4858 */;
                4631: data_o = 32'h00000000 /* 0x485c */;
                4632: data_o = 32'h00000000 /* 0x4860 */;
                4633: data_o = 32'h00000000 /* 0x4864 */;
                4634: data_o = 32'h00000000 /* 0x4868 */;
                4635: data_o = 32'h00000000 /* 0x486c */;
                4636: data_o = 32'h00000000 /* 0x4870 */;
                4637: data_o = 32'h00000000 /* 0x4874 */;
                4638: data_o = 32'h00000000 /* 0x4878 */;
                4639: data_o = 32'h00000000 /* 0x487c */;
                4640: data_o = 32'h00000000 /* 0x4880 */;
                4641: data_o = 32'h00000000 /* 0x4884 */;
                4642: data_o = 32'h00000000 /* 0x4888 */;
                4643: data_o = 32'h00000000 /* 0x488c */;
                4644: data_o = 32'h00000000 /* 0x4890 */;
                4645: data_o = 32'h00000000 /* 0x4894 */;
                4646: data_o = 32'h00000000 /* 0x4898 */;
                4647: data_o = 32'h00000000 /* 0x489c */;
                4648: data_o = 32'h00000000 /* 0x48a0 */;
                4649: data_o = 32'h00000000 /* 0x48a4 */;
                4650: data_o = 32'h00000000 /* 0x48a8 */;
                4651: data_o = 32'h00000000 /* 0x48ac */;
                4652: data_o = 32'h00000000 /* 0x48b0 */;
                4653: data_o = 32'h00000000 /* 0x48b4 */;
                4654: data_o = 32'h00000000 /* 0x48b8 */;
                4655: data_o = 32'h00000000 /* 0x48bc */;
                4656: data_o = 32'h00000000 /* 0x48c0 */;
                4657: data_o = 32'h00000000 /* 0x48c4 */;
                4658: data_o = 32'h00000000 /* 0x48c8 */;
                4659: data_o = 32'h00000000 /* 0x48cc */;
                4660: data_o = 32'h00000000 /* 0x48d0 */;
                4661: data_o = 32'h00000000 /* 0x48d4 */;
                4662: data_o = 32'h00000000 /* 0x48d8 */;
                4663: data_o = 32'h00000000 /* 0x48dc */;
                4664: data_o = 32'h00000000 /* 0x48e0 */;
                4665: data_o = 32'h00000000 /* 0x48e4 */;
                4666: data_o = 32'h00000000 /* 0x48e8 */;
                4667: data_o = 32'h00000000 /* 0x48ec */;
                4668: data_o = 32'h00000000 /* 0x48f0 */;
                4669: data_o = 32'h00000000 /* 0x48f4 */;
                4670: data_o = 32'h00000000 /* 0x48f8 */;
                4671: data_o = 32'h00000000 /* 0x48fc */;
                4672: data_o = 32'h00000000 /* 0x4900 */;
                4673: data_o = 32'h00000000 /* 0x4904 */;
                4674: data_o = 32'h00000000 /* 0x4908 */;
                4675: data_o = 32'h00000000 /* 0x490c */;
                4676: data_o = 32'h00000000 /* 0x4910 */;
                4677: data_o = 32'h00000000 /* 0x4914 */;
                4678: data_o = 32'h00000000 /* 0x4918 */;
                4679: data_o = 32'h00000000 /* 0x491c */;
                4680: data_o = 32'h00000000 /* 0x4920 */;
                4681: data_o = 32'h00000000 /* 0x4924 */;
                4682: data_o = 32'h00000000 /* 0x4928 */;
                4683: data_o = 32'h00000000 /* 0x492c */;
                4684: data_o = 32'h00000000 /* 0x4930 */;
                4685: data_o = 32'h00000000 /* 0x4934 */;
                4686: data_o = 32'h00000000 /* 0x4938 */;
                4687: data_o = 32'h00000000 /* 0x493c */;
                4688: data_o = 32'h00000000 /* 0x4940 */;
                4689: data_o = 32'h00000000 /* 0x4944 */;
                4690: data_o = 32'h00000000 /* 0x4948 */;
                4691: data_o = 32'h00000000 /* 0x494c */;
                4692: data_o = 32'h00000000 /* 0x4950 */;
                4693: data_o = 32'h00000000 /* 0x4954 */;
                4694: data_o = 32'h00000000 /* 0x4958 */;
                4695: data_o = 32'h00000000 /* 0x495c */;
                4696: data_o = 32'h00000000 /* 0x4960 */;
                4697: data_o = 32'h00000000 /* 0x4964 */;
                4698: data_o = 32'h00000000 /* 0x4968 */;
                4699: data_o = 32'h00000000 /* 0x496c */;
                4700: data_o = 32'h00000000 /* 0x4970 */;
                4701: data_o = 32'h00000000 /* 0x4974 */;
                4702: data_o = 32'h00000000 /* 0x4978 */;
                4703: data_o = 32'h00000000 /* 0x497c */;
                4704: data_o = 32'h00000000 /* 0x4980 */;
                4705: data_o = 32'h00000000 /* 0x4984 */;
                4706: data_o = 32'h00000000 /* 0x4988 */;
                4707: data_o = 32'h00000000 /* 0x498c */;
                4708: data_o = 32'h00000000 /* 0x4990 */;
                4709: data_o = 32'h00000000 /* 0x4994 */;
                4710: data_o = 32'h00000000 /* 0x4998 */;
                4711: data_o = 32'h00000000 /* 0x499c */;
                4712: data_o = 32'h00000000 /* 0x49a0 */;
                4713: data_o = 32'h00000000 /* 0x49a4 */;
                4714: data_o = 32'h00000000 /* 0x49a8 */;
                4715: data_o = 32'h00000000 /* 0x49ac */;
                4716: data_o = 32'h00000000 /* 0x49b0 */;
                4717: data_o = 32'h00000000 /* 0x49b4 */;
                4718: data_o = 32'h00000000 /* 0x49b8 */;
                4719: data_o = 32'h00000000 /* 0x49bc */;
                4720: data_o = 32'h00000000 /* 0x49c0 */;
                4721: data_o = 32'h00000000 /* 0x49c4 */;
                4722: data_o = 32'h00000000 /* 0x49c8 */;
                4723: data_o = 32'h00000000 /* 0x49cc */;
                4724: data_o = 32'h00000000 /* 0x49d0 */;
                4725: data_o = 32'h00000000 /* 0x49d4 */;
                4726: data_o = 32'h00000000 /* 0x49d8 */;
                4727: data_o = 32'h00000000 /* 0x49dc */;
                4728: data_o = 32'h00000000 /* 0x49e0 */;
                4729: data_o = 32'h00000000 /* 0x49e4 */;
                4730: data_o = 32'h00000000 /* 0x49e8 */;
                4731: data_o = 32'h00000000 /* 0x49ec */;
                4732: data_o = 32'h00000000 /* 0x49f0 */;
                4733: data_o = 32'h00000000 /* 0x49f4 */;
                4734: data_o = 32'h00000000 /* 0x49f8 */;
                4735: data_o = 32'h00000000 /* 0x49fc */;
                4736: data_o = 32'h00000000 /* 0x4a00 */;
                4737: data_o = 32'h00000000 /* 0x4a04 */;
                4738: data_o = 32'h00000000 /* 0x4a08 */;
                4739: data_o = 32'h00000000 /* 0x4a0c */;
                4740: data_o = 32'h00000000 /* 0x4a10 */;
                4741: data_o = 32'h00000000 /* 0x4a14 */;
                4742: data_o = 32'h00000000 /* 0x4a18 */;
                4743: data_o = 32'h00000000 /* 0x4a1c */;
                4744: data_o = 32'h00000000 /* 0x4a20 */;
                4745: data_o = 32'h00000000 /* 0x4a24 */;
                4746: data_o = 32'h00000000 /* 0x4a28 */;
                4747: data_o = 32'h00000000 /* 0x4a2c */;
                4748: data_o = 32'h00000000 /* 0x4a30 */;
                4749: data_o = 32'h00000000 /* 0x4a34 */;
                4750: data_o = 32'h00000000 /* 0x4a38 */;
                4751: data_o = 32'h00000000 /* 0x4a3c */;
                4752: data_o = 32'h00000000 /* 0x4a40 */;
                4753: data_o = 32'h00000000 /* 0x4a44 */;
                4754: data_o = 32'h00000000 /* 0x4a48 */;
                4755: data_o = 32'h00000000 /* 0x4a4c */;
                4756: data_o = 32'h00000000 /* 0x4a50 */;
                4757: data_o = 32'h00000000 /* 0x4a54 */;
                4758: data_o = 32'h00000000 /* 0x4a58 */;
                4759: data_o = 32'h00000000 /* 0x4a5c */;
                4760: data_o = 32'h00000000 /* 0x4a60 */;
                4761: data_o = 32'h00000000 /* 0x4a64 */;
                4762: data_o = 32'h00000000 /* 0x4a68 */;
                4763: data_o = 32'h00000000 /* 0x4a6c */;
                4764: data_o = 32'h00000000 /* 0x4a70 */;
                4765: data_o = 32'h00000000 /* 0x4a74 */;
                4766: data_o = 32'h00000000 /* 0x4a78 */;
                4767: data_o = 32'h00000000 /* 0x4a7c */;
                4768: data_o = 32'h00000000 /* 0x4a80 */;
                4769: data_o = 32'h00000000 /* 0x4a84 */;
                4770: data_o = 32'h00000000 /* 0x4a88 */;
                4771: data_o = 32'h00000000 /* 0x4a8c */;
                4772: data_o = 32'h00000000 /* 0x4a90 */;
                4773: data_o = 32'h00000000 /* 0x4a94 */;
                4774: data_o = 32'h00000000 /* 0x4a98 */;
                4775: data_o = 32'h00000000 /* 0x4a9c */;
                4776: data_o = 32'h00000000 /* 0x4aa0 */;
                4777: data_o = 32'h00000000 /* 0x4aa4 */;
                4778: data_o = 32'h00000000 /* 0x4aa8 */;
                4779: data_o = 32'h00000000 /* 0x4aac */;
                4780: data_o = 32'h00000000 /* 0x4ab0 */;
                4781: data_o = 32'h00000000 /* 0x4ab4 */;
                4782: data_o = 32'h00000000 /* 0x4ab8 */;
                4783: data_o = 32'h00000000 /* 0x4abc */;
                4784: data_o = 32'h00000000 /* 0x4ac0 */;
                4785: data_o = 32'h00000000 /* 0x4ac4 */;
                4786: data_o = 32'h00000000 /* 0x4ac8 */;
                4787: data_o = 32'h00000000 /* 0x4acc */;
                4788: data_o = 32'h00000000 /* 0x4ad0 */;
                4789: data_o = 32'h00000000 /* 0x4ad4 */;
                4790: data_o = 32'h00000000 /* 0x4ad8 */;
                4791: data_o = 32'h00000000 /* 0x4adc */;
                4792: data_o = 32'h00000000 /* 0x4ae0 */;
                4793: data_o = 32'h00000000 /* 0x4ae4 */;
                4794: data_o = 32'h00000000 /* 0x4ae8 */;
                4795: data_o = 32'h00000000 /* 0x4aec */;
                4796: data_o = 32'h00000000 /* 0x4af0 */;
                4797: data_o = 32'h00000000 /* 0x4af4 */;
                4798: data_o = 32'h00000000 /* 0x4af8 */;
                4799: data_o = 32'h00000000 /* 0x4afc */;
                4800: data_o = 32'h00000000 /* 0x4b00 */;
                4801: data_o = 32'h00000000 /* 0x4b04 */;
                4802: data_o = 32'h00000000 /* 0x4b08 */;
                4803: data_o = 32'h00000000 /* 0x4b0c */;
                4804: data_o = 32'h00000000 /* 0x4b10 */;
                4805: data_o = 32'h00000000 /* 0x4b14 */;
                4806: data_o = 32'h00000000 /* 0x4b18 */;
                4807: data_o = 32'h00000000 /* 0x4b1c */;
                4808: data_o = 32'h00000000 /* 0x4b20 */;
                4809: data_o = 32'h00000000 /* 0x4b24 */;
                4810: data_o = 32'h00000000 /* 0x4b28 */;
                4811: data_o = 32'h00000000 /* 0x4b2c */;
                4812: data_o = 32'h00000000 /* 0x4b30 */;
                4813: data_o = 32'h00000000 /* 0x4b34 */;
                4814: data_o = 32'h00000000 /* 0x4b38 */;
                4815: data_o = 32'h00000000 /* 0x4b3c */;
                4816: data_o = 32'h00000000 /* 0x4b40 */;
                4817: data_o = 32'h00000000 /* 0x4b44 */;
                4818: data_o = 32'h00000000 /* 0x4b48 */;
                4819: data_o = 32'h00000000 /* 0x4b4c */;
                4820: data_o = 32'h00000000 /* 0x4b50 */;
                4821: data_o = 32'h00000000 /* 0x4b54 */;
                4822: data_o = 32'h00000000 /* 0x4b58 */;
                4823: data_o = 32'h00000000 /* 0x4b5c */;
                4824: data_o = 32'h00000000 /* 0x4b60 */;
                4825: data_o = 32'h00000000 /* 0x4b64 */;
                4826: data_o = 32'h00000000 /* 0x4b68 */;
                4827: data_o = 32'h00000000 /* 0x4b6c */;
                4828: data_o = 32'h00000000 /* 0x4b70 */;
                4829: data_o = 32'h00000000 /* 0x4b74 */;
                4830: data_o = 32'h00000000 /* 0x4b78 */;
                4831: data_o = 32'h00000000 /* 0x4b7c */;
                4832: data_o = 32'h00000000 /* 0x4b80 */;
                4833: data_o = 32'h00000000 /* 0x4b84 */;
                4834: data_o = 32'h00000000 /* 0x4b88 */;
                4835: data_o = 32'h00000000 /* 0x4b8c */;
                4836: data_o = 32'h00000000 /* 0x4b90 */;
                4837: data_o = 32'h00000000 /* 0x4b94 */;
                4838: data_o = 32'h00000000 /* 0x4b98 */;
                4839: data_o = 32'h00000000 /* 0x4b9c */;
                4840: data_o = 32'h00000000 /* 0x4ba0 */;
                4841: data_o = 32'h00000000 /* 0x4ba4 */;
                4842: data_o = 32'h00000000 /* 0x4ba8 */;
                4843: data_o = 32'h00000000 /* 0x4bac */;
                4844: data_o = 32'h00000000 /* 0x4bb0 */;
                4845: data_o = 32'h00000000 /* 0x4bb4 */;
                4846: data_o = 32'h00000000 /* 0x4bb8 */;
                4847: data_o = 32'h00000000 /* 0x4bbc */;
                4848: data_o = 32'h00000000 /* 0x4bc0 */;
                4849: data_o = 32'h00000000 /* 0x4bc4 */;
                4850: data_o = 32'h00000000 /* 0x4bc8 */;
                4851: data_o = 32'h00000000 /* 0x4bcc */;
                4852: data_o = 32'h00000000 /* 0x4bd0 */;
                4853: data_o = 32'h00000000 /* 0x4bd4 */;
                4854: data_o = 32'h00000000 /* 0x4bd8 */;
                4855: data_o = 32'h00000000 /* 0x4bdc */;
                4856: data_o = 32'h00000000 /* 0x4be0 */;
                4857: data_o = 32'h00000000 /* 0x4be4 */;
                4858: data_o = 32'h00000000 /* 0x4be8 */;
                4859: data_o = 32'h00000000 /* 0x4bec */;
                4860: data_o = 32'h00000000 /* 0x4bf0 */;
                4861: data_o = 32'h00000000 /* 0x4bf4 */;
                4862: data_o = 32'h00000000 /* 0x4bf8 */;
                4863: data_o = 32'h00000000 /* 0x4bfc */;
                4864: data_o = 32'h00000000 /* 0x4c00 */;
                4865: data_o = 32'h00000000 /* 0x4c04 */;
                4866: data_o = 32'h00000000 /* 0x4c08 */;
                4867: data_o = 32'h00000000 /* 0x4c0c */;
                4868: data_o = 32'h00000000 /* 0x4c10 */;
                4869: data_o = 32'h00000000 /* 0x4c14 */;
                4870: data_o = 32'h00000000 /* 0x4c18 */;
                4871: data_o = 32'h00000000 /* 0x4c1c */;
                4872: data_o = 32'h00000000 /* 0x4c20 */;
                4873: data_o = 32'h00000000 /* 0x4c24 */;
                4874: data_o = 32'h00000000 /* 0x4c28 */;
                4875: data_o = 32'h00000000 /* 0x4c2c */;
                4876: data_o = 32'h00000000 /* 0x4c30 */;
                4877: data_o = 32'h00000000 /* 0x4c34 */;
                4878: data_o = 32'h00000000 /* 0x4c38 */;
                4879: data_o = 32'h00000000 /* 0x4c3c */;
                4880: data_o = 32'h00000000 /* 0x4c40 */;
                4881: data_o = 32'h00000000 /* 0x4c44 */;
                4882: data_o = 32'h00000000 /* 0x4c48 */;
                4883: data_o = 32'h00000000 /* 0x4c4c */;
                4884: data_o = 32'h00000000 /* 0x4c50 */;
                4885: data_o = 32'h00000000 /* 0x4c54 */;
                4886: data_o = 32'h00000000 /* 0x4c58 */;
                4887: data_o = 32'h00000000 /* 0x4c5c */;
                4888: data_o = 32'h00000000 /* 0x4c60 */;
                4889: data_o = 32'h00000000 /* 0x4c64 */;
                4890: data_o = 32'h00000000 /* 0x4c68 */;
                4891: data_o = 32'h00000000 /* 0x4c6c */;
                4892: data_o = 32'h00000000 /* 0x4c70 */;
                4893: data_o = 32'h00000000 /* 0x4c74 */;
                4894: data_o = 32'h00000000 /* 0x4c78 */;
                4895: data_o = 32'h00000000 /* 0x4c7c */;
                4896: data_o = 32'h00000000 /* 0x4c80 */;
                4897: data_o = 32'h00000000 /* 0x4c84 */;
                4898: data_o = 32'h00000000 /* 0x4c88 */;
                4899: data_o = 32'h00000000 /* 0x4c8c */;
                4900: data_o = 32'h00000000 /* 0x4c90 */;
                4901: data_o = 32'h00000000 /* 0x4c94 */;
                4902: data_o = 32'h00000000 /* 0x4c98 */;
                4903: data_o = 32'h00000000 /* 0x4c9c */;
                4904: data_o = 32'h00000000 /* 0x4ca0 */;
                4905: data_o = 32'h00000000 /* 0x4ca4 */;
                4906: data_o = 32'h00000000 /* 0x4ca8 */;
                4907: data_o = 32'h00000000 /* 0x4cac */;
                4908: data_o = 32'h00000000 /* 0x4cb0 */;
                4909: data_o = 32'h00000000 /* 0x4cb4 */;
                4910: data_o = 32'h00000000 /* 0x4cb8 */;
                4911: data_o = 32'h00000000 /* 0x4cbc */;
                4912: data_o = 32'h00000000 /* 0x4cc0 */;
                4913: data_o = 32'h00000000 /* 0x4cc4 */;
                4914: data_o = 32'h00000000 /* 0x4cc8 */;
                4915: data_o = 32'h00000000 /* 0x4ccc */;
                4916: data_o = 32'h00000000 /* 0x4cd0 */;
                4917: data_o = 32'h00000000 /* 0x4cd4 */;
                4918: data_o = 32'h00000000 /* 0x4cd8 */;
                4919: data_o = 32'h00000000 /* 0x4cdc */;
                4920: data_o = 32'h00000000 /* 0x4ce0 */;
                4921: data_o = 32'h00000000 /* 0x4ce4 */;
                4922: data_o = 32'h00000000 /* 0x4ce8 */;
                4923: data_o = 32'h00000000 /* 0x4cec */;
                4924: data_o = 32'h00000000 /* 0x4cf0 */;
                4925: data_o = 32'h00000000 /* 0x4cf4 */;
                4926: data_o = 32'h00000000 /* 0x4cf8 */;
                4927: data_o = 32'h00000000 /* 0x4cfc */;
                4928: data_o = 32'h00000000 /* 0x4d00 */;
                4929: data_o = 32'h00000000 /* 0x4d04 */;
                4930: data_o = 32'h00000000 /* 0x4d08 */;
                4931: data_o = 32'h00000000 /* 0x4d0c */;
                4932: data_o = 32'h00000000 /* 0x4d10 */;
                4933: data_o = 32'h00000000 /* 0x4d14 */;
                4934: data_o = 32'h00000000 /* 0x4d18 */;
                4935: data_o = 32'h00000000 /* 0x4d1c */;
                4936: data_o = 32'h00000000 /* 0x4d20 */;
                4937: data_o = 32'h00000000 /* 0x4d24 */;
                4938: data_o = 32'h00000000 /* 0x4d28 */;
                4939: data_o = 32'h00000000 /* 0x4d2c */;
                4940: data_o = 32'h00000000 /* 0x4d30 */;
                4941: data_o = 32'h00000000 /* 0x4d34 */;
                4942: data_o = 32'h00000000 /* 0x4d38 */;
                4943: data_o = 32'h00000000 /* 0x4d3c */;
                4944: data_o = 32'h00000000 /* 0x4d40 */;
                4945: data_o = 32'h00000000 /* 0x4d44 */;
                4946: data_o = 32'h00000000 /* 0x4d48 */;
                4947: data_o = 32'h00000000 /* 0x4d4c */;
                4948: data_o = 32'h00000000 /* 0x4d50 */;
                4949: data_o = 32'h00000000 /* 0x4d54 */;
                4950: data_o = 32'h00000000 /* 0x4d58 */;
                4951: data_o = 32'h00000000 /* 0x4d5c */;
                4952: data_o = 32'h00000000 /* 0x4d60 */;
                4953: data_o = 32'h00000000 /* 0x4d64 */;
                4954: data_o = 32'h00000000 /* 0x4d68 */;
                4955: data_o = 32'h00000000 /* 0x4d6c */;
                4956: data_o = 32'h00000000 /* 0x4d70 */;
                4957: data_o = 32'h00000000 /* 0x4d74 */;
                4958: data_o = 32'h00000000 /* 0x4d78 */;
                4959: data_o = 32'h00000000 /* 0x4d7c */;
                4960: data_o = 32'h00000000 /* 0x4d80 */;
                4961: data_o = 32'h00000000 /* 0x4d84 */;
                4962: data_o = 32'h00000000 /* 0x4d88 */;
                4963: data_o = 32'h00000000 /* 0x4d8c */;
                4964: data_o = 32'h00000000 /* 0x4d90 */;
                4965: data_o = 32'h00000000 /* 0x4d94 */;
                4966: data_o = 32'h00000000 /* 0x4d98 */;
                4967: data_o = 32'h00000000 /* 0x4d9c */;
                4968: data_o = 32'h00000000 /* 0x4da0 */;
                4969: data_o = 32'h00000000 /* 0x4da4 */;
                4970: data_o = 32'h00000000 /* 0x4da8 */;
                4971: data_o = 32'h00000000 /* 0x4dac */;
                4972: data_o = 32'h00000000 /* 0x4db0 */;
                4973: data_o = 32'h00000000 /* 0x4db4 */;
                4974: data_o = 32'h00000000 /* 0x4db8 */;
                4975: data_o = 32'h00000000 /* 0x4dbc */;
                4976: data_o = 32'h00000000 /* 0x4dc0 */;
                4977: data_o = 32'h00000000 /* 0x4dc4 */;
                4978: data_o = 32'h00000000 /* 0x4dc8 */;
                4979: data_o = 32'h00000000 /* 0x4dcc */;
                4980: data_o = 32'h00000000 /* 0x4dd0 */;
                4981: data_o = 32'h00000000 /* 0x4dd4 */;
                4982: data_o = 32'h00000000 /* 0x4dd8 */;
                4983: data_o = 32'h00000000 /* 0x4ddc */;
                4984: data_o = 32'h00000000 /* 0x4de0 */;
                4985: data_o = 32'h00000000 /* 0x4de4 */;
                4986: data_o = 32'h00000000 /* 0x4de8 */;
                4987: data_o = 32'h00000000 /* 0x4dec */;
                4988: data_o = 32'h00000000 /* 0x4df0 */;
                4989: data_o = 32'h00000000 /* 0x4df4 */;
                4990: data_o = 32'h00000000 /* 0x4df8 */;
                4991: data_o = 32'h00000000 /* 0x4dfc */;
                4992: data_o = 32'h00000000 /* 0x4e00 */;
                4993: data_o = 32'h00000000 /* 0x4e04 */;
                4994: data_o = 32'h00000000 /* 0x4e08 */;
                4995: data_o = 32'h00000000 /* 0x4e0c */;
                4996: data_o = 32'h00000000 /* 0x4e10 */;
                4997: data_o = 32'h00000000 /* 0x4e14 */;
                4998: data_o = 32'h00000000 /* 0x4e18 */;
                4999: data_o = 32'h00000000 /* 0x4e1c */;
                5000: data_o = 32'h00000000 /* 0x4e20 */;
                5001: data_o = 32'h00000000 /* 0x4e24 */;
                5002: data_o = 32'h00000000 /* 0x4e28 */;
                5003: data_o = 32'h00000000 /* 0x4e2c */;
                5004: data_o = 32'h00000000 /* 0x4e30 */;
                5005: data_o = 32'h00000000 /* 0x4e34 */;
                5006: data_o = 32'h00000000 /* 0x4e38 */;
                5007: data_o = 32'h00000000 /* 0x4e3c */;
                5008: data_o = 32'h00000000 /* 0x4e40 */;
                5009: data_o = 32'h00000000 /* 0x4e44 */;
                5010: data_o = 32'h00000000 /* 0x4e48 */;
                5011: data_o = 32'h00000000 /* 0x4e4c */;
                5012: data_o = 32'h00000000 /* 0x4e50 */;
                5013: data_o = 32'h00000000 /* 0x4e54 */;
                5014: data_o = 32'h00000000 /* 0x4e58 */;
                5015: data_o = 32'h00000000 /* 0x4e5c */;
                5016: data_o = 32'h00000000 /* 0x4e60 */;
                5017: data_o = 32'h00000000 /* 0x4e64 */;
                5018: data_o = 32'h00000000 /* 0x4e68 */;
                5019: data_o = 32'h00000000 /* 0x4e6c */;
                5020: data_o = 32'h00000000 /* 0x4e70 */;
                5021: data_o = 32'h00000000 /* 0x4e74 */;
                5022: data_o = 32'h00000000 /* 0x4e78 */;
                5023: data_o = 32'h00000000 /* 0x4e7c */;
                5024: data_o = 32'h00000000 /* 0x4e80 */;
                5025: data_o = 32'h00000000 /* 0x4e84 */;
                5026: data_o = 32'h00000000 /* 0x4e88 */;
                5027: data_o = 32'h00000000 /* 0x4e8c */;
                5028: data_o = 32'h00000000 /* 0x4e90 */;
                5029: data_o = 32'h00000000 /* 0x4e94 */;
                5030: data_o = 32'h00000000 /* 0x4e98 */;
                5031: data_o = 32'h00000000 /* 0x4e9c */;
                5032: data_o = 32'h00000000 /* 0x4ea0 */;
                5033: data_o = 32'h00000000 /* 0x4ea4 */;
                5034: data_o = 32'h00000000 /* 0x4ea8 */;
                5035: data_o = 32'h00000000 /* 0x4eac */;
                5036: data_o = 32'h00000000 /* 0x4eb0 */;
                5037: data_o = 32'h00000000 /* 0x4eb4 */;
                5038: data_o = 32'h00000000 /* 0x4eb8 */;
                5039: data_o = 32'h00000000 /* 0x4ebc */;
                5040: data_o = 32'h00000000 /* 0x4ec0 */;
                5041: data_o = 32'h00000000 /* 0x4ec4 */;
                5042: data_o = 32'h00000000 /* 0x4ec8 */;
                5043: data_o = 32'h00000000 /* 0x4ecc */;
                5044: data_o = 32'h00000000 /* 0x4ed0 */;
                5045: data_o = 32'h00000000 /* 0x4ed4 */;
                5046: data_o = 32'h00000000 /* 0x4ed8 */;
                5047: data_o = 32'h00000000 /* 0x4edc */;
                5048: data_o = 32'h00000000 /* 0x4ee0 */;
                5049: data_o = 32'h00000000 /* 0x4ee4 */;
                5050: data_o = 32'h00000000 /* 0x4ee8 */;
                5051: data_o = 32'h00000000 /* 0x4eec */;
                5052: data_o = 32'h00000000 /* 0x4ef0 */;
                5053: data_o = 32'h00000000 /* 0x4ef4 */;
                5054: data_o = 32'h00000000 /* 0x4ef8 */;
                5055: data_o = 32'h00000000 /* 0x4efc */;
                5056: data_o = 32'h00000000 /* 0x4f00 */;
                5057: data_o = 32'h00000000 /* 0x4f04 */;
                5058: data_o = 32'h00000000 /* 0x4f08 */;
                5059: data_o = 32'h00000000 /* 0x4f0c */;
                5060: data_o = 32'h00000000 /* 0x4f10 */;
                5061: data_o = 32'h00000000 /* 0x4f14 */;
                5062: data_o = 32'h00000000 /* 0x4f18 */;
                5063: data_o = 32'h00000000 /* 0x4f1c */;
                5064: data_o = 32'h00000000 /* 0x4f20 */;
                5065: data_o = 32'h00000000 /* 0x4f24 */;
                5066: data_o = 32'h00000000 /* 0x4f28 */;
                5067: data_o = 32'h00000000 /* 0x4f2c */;
                5068: data_o = 32'h00000000 /* 0x4f30 */;
                5069: data_o = 32'h00000000 /* 0x4f34 */;
                5070: data_o = 32'h00000000 /* 0x4f38 */;
                5071: data_o = 32'h00000000 /* 0x4f3c */;
                5072: data_o = 32'h00000000 /* 0x4f40 */;
                5073: data_o = 32'h00000000 /* 0x4f44 */;
                5074: data_o = 32'h00000000 /* 0x4f48 */;
                5075: data_o = 32'h00000000 /* 0x4f4c */;
                5076: data_o = 32'h00000000 /* 0x4f50 */;
                5077: data_o = 32'h00000000 /* 0x4f54 */;
                5078: data_o = 32'h00000000 /* 0x4f58 */;
                5079: data_o = 32'h00000000 /* 0x4f5c */;
                5080: data_o = 32'h00000000 /* 0x4f60 */;
                5081: data_o = 32'h00000000 /* 0x4f64 */;
                5082: data_o = 32'h00000000 /* 0x4f68 */;
                5083: data_o = 32'h00000000 /* 0x4f6c */;
                5084: data_o = 32'h00000000 /* 0x4f70 */;
                5085: data_o = 32'h00000000 /* 0x4f74 */;
                5086: data_o = 32'h00000000 /* 0x4f78 */;
                5087: data_o = 32'h00000000 /* 0x4f7c */;
                5088: data_o = 32'h00000000 /* 0x4f80 */;
                5089: data_o = 32'h00000000 /* 0x4f84 */;
                5090: data_o = 32'h00000000 /* 0x4f88 */;
                5091: data_o = 32'h00000000 /* 0x4f8c */;
                5092: data_o = 32'h00000000 /* 0x4f90 */;
                5093: data_o = 32'h00000000 /* 0x4f94 */;
                5094: data_o = 32'h00000000 /* 0x4f98 */;
                5095: data_o = 32'h00000000 /* 0x4f9c */;
                5096: data_o = 32'h00000000 /* 0x4fa0 */;
                5097: data_o = 32'h00000000 /* 0x4fa4 */;
                5098: data_o = 32'h00000000 /* 0x4fa8 */;
                5099: data_o = 32'h00000000 /* 0x4fac */;
                5100: data_o = 32'h00000000 /* 0x4fb0 */;
                5101: data_o = 32'h00000000 /* 0x4fb4 */;
                5102: data_o = 32'h00000000 /* 0x4fb8 */;
                5103: data_o = 32'h00000000 /* 0x4fbc */;
                5104: data_o = 32'h00000000 /* 0x4fc0 */;
                5105: data_o = 32'h00000000 /* 0x4fc4 */;
                5106: data_o = 32'h00000000 /* 0x4fc8 */;
                5107: data_o = 32'h00000000 /* 0x4fcc */;
                5108: data_o = 32'h00000000 /* 0x4fd0 */;
                5109: data_o = 32'h00000000 /* 0x4fd4 */;
                5110: data_o = 32'h00000000 /* 0x4fd8 */;
                5111: data_o = 32'h00000000 /* 0x4fdc */;
                5112: data_o = 32'h00000000 /* 0x4fe0 */;
                5113: data_o = 32'h00000000 /* 0x4fe4 */;
                5114: data_o = 32'h00000000 /* 0x4fe8 */;
                5115: data_o = 32'h00000000 /* 0x4fec */;
                5116: data_o = 32'h00000000 /* 0x4ff0 */;
                5117: data_o = 32'h00000000 /* 0x4ff4 */;
                5118: data_o = 32'h00000000 /* 0x4ff8 */;
                5119: data_o = 32'h00000000 /* 0x4ffc */;
                5120: data_o = 32'h00000000 /* 0x5000 */;
                5121: data_o = 32'h00000000 /* 0x5004 */;
                5122: data_o = 32'h00000000 /* 0x5008 */;
                5123: data_o = 32'h00000000 /* 0x500c */;
                5124: data_o = 32'h00000000 /* 0x5010 */;
                5125: data_o = 32'h00000000 /* 0x5014 */;
                5126: data_o = 32'h00000000 /* 0x5018 */;
                5127: data_o = 32'h00000000 /* 0x501c */;
                5128: data_o = 32'h00000000 /* 0x5020 */;
                5129: data_o = 32'h00000000 /* 0x5024 */;
                5130: data_o = 32'h00000000 /* 0x5028 */;
                5131: data_o = 32'h00000000 /* 0x502c */;
                5132: data_o = 32'h00000000 /* 0x5030 */;
                5133: data_o = 32'h00000000 /* 0x5034 */;
                5134: data_o = 32'h00000000 /* 0x5038 */;
                5135: data_o = 32'h00000000 /* 0x503c */;
                5136: data_o = 32'h00000000 /* 0x5040 */;
                5137: data_o = 32'h00000000 /* 0x5044 */;
                5138: data_o = 32'h00000000 /* 0x5048 */;
                5139: data_o = 32'h00000000 /* 0x504c */;
                5140: data_o = 32'h00000000 /* 0x5050 */;
                5141: data_o = 32'h00000000 /* 0x5054 */;
                5142: data_o = 32'h00000000 /* 0x5058 */;
                5143: data_o = 32'h00000000 /* 0x505c */;
                5144: data_o = 32'h00000000 /* 0x5060 */;
                5145: data_o = 32'h00000000 /* 0x5064 */;
                5146: data_o = 32'h00000000 /* 0x5068 */;
                5147: data_o = 32'h00000000 /* 0x506c */;
                5148: data_o = 32'h00000000 /* 0x5070 */;
                5149: data_o = 32'h00000000 /* 0x5074 */;
                5150: data_o = 32'h00000000 /* 0x5078 */;
                5151: data_o = 32'h00000000 /* 0x507c */;
                5152: data_o = 32'h00000000 /* 0x5080 */;
                5153: data_o = 32'h00000000 /* 0x5084 */;
                5154: data_o = 32'h00000000 /* 0x5088 */;
                5155: data_o = 32'h00000000 /* 0x508c */;
                5156: data_o = 32'h00000000 /* 0x5090 */;
                5157: data_o = 32'h00000000 /* 0x5094 */;
                5158: data_o = 32'h00000000 /* 0x5098 */;
                5159: data_o = 32'h00000000 /* 0x509c */;
                5160: data_o = 32'h00000000 /* 0x50a0 */;
                5161: data_o = 32'h00000000 /* 0x50a4 */;
                5162: data_o = 32'h00000000 /* 0x50a8 */;
                5163: data_o = 32'h00000000 /* 0x50ac */;
                5164: data_o = 32'h00000000 /* 0x50b0 */;
                5165: data_o = 32'h00000000 /* 0x50b4 */;
                5166: data_o = 32'h00000000 /* 0x50b8 */;
                5167: data_o = 32'h00000000 /* 0x50bc */;
                5168: data_o = 32'h00000000 /* 0x50c0 */;
                5169: data_o = 32'h00000000 /* 0x50c4 */;
                5170: data_o = 32'h00000000 /* 0x50c8 */;
                5171: data_o = 32'h00000000 /* 0x50cc */;
                5172: data_o = 32'h00000000 /* 0x50d0 */;
                5173: data_o = 32'h00000000 /* 0x50d4 */;
                5174: data_o = 32'h00000000 /* 0x50d8 */;
                5175: data_o = 32'h00000000 /* 0x50dc */;
                5176: data_o = 32'h00000000 /* 0x50e0 */;
                5177: data_o = 32'h00000000 /* 0x50e4 */;
                5178: data_o = 32'h00000000 /* 0x50e8 */;
                5179: data_o = 32'h00000000 /* 0x50ec */;
                5180: data_o = 32'h00000000 /* 0x50f0 */;
                5181: data_o = 32'h00000000 /* 0x50f4 */;
                5182: data_o = 32'h00000000 /* 0x50f8 */;
                5183: data_o = 32'h00000000 /* 0x50fc */;
                5184: data_o = 32'h00000000 /* 0x5100 */;
                5185: data_o = 32'h00000000 /* 0x5104 */;
                5186: data_o = 32'h00000000 /* 0x5108 */;
                5187: data_o = 32'h00000000 /* 0x510c */;
                5188: data_o = 32'h00000000 /* 0x5110 */;
                5189: data_o = 32'h00000000 /* 0x5114 */;
                5190: data_o = 32'h00000000 /* 0x5118 */;
                5191: data_o = 32'h00000000 /* 0x511c */;
                5192: data_o = 32'h00000000 /* 0x5120 */;
                5193: data_o = 32'h00000000 /* 0x5124 */;
                5194: data_o = 32'h00000000 /* 0x5128 */;
                5195: data_o = 32'h00000000 /* 0x512c */;
                5196: data_o = 32'h00000000 /* 0x5130 */;
                5197: data_o = 32'h00000000 /* 0x5134 */;
                5198: data_o = 32'h00000000 /* 0x5138 */;
                5199: data_o = 32'h00000000 /* 0x513c */;
                5200: data_o = 32'h00000000 /* 0x5140 */;
                5201: data_o = 32'h00000000 /* 0x5144 */;
                5202: data_o = 32'h00000000 /* 0x5148 */;
                5203: data_o = 32'h00000000 /* 0x514c */;
                5204: data_o = 32'h00000000 /* 0x5150 */;
                5205: data_o = 32'h00000000 /* 0x5154 */;
                5206: data_o = 32'h00000000 /* 0x5158 */;
                5207: data_o = 32'h00000000 /* 0x515c */;
                5208: data_o = 32'h00000000 /* 0x5160 */;
                5209: data_o = 32'h00000000 /* 0x5164 */;
                5210: data_o = 32'h00000000 /* 0x5168 */;
                5211: data_o = 32'h00000000 /* 0x516c */;
                5212: data_o = 32'h00000000 /* 0x5170 */;
                5213: data_o = 32'h00000000 /* 0x5174 */;
                5214: data_o = 32'h00000000 /* 0x5178 */;
                5215: data_o = 32'h00000000 /* 0x517c */;
                5216: data_o = 32'h00000000 /* 0x5180 */;
                5217: data_o = 32'h00000000 /* 0x5184 */;
                5218: data_o = 32'h00000000 /* 0x5188 */;
                5219: data_o = 32'h00000000 /* 0x518c */;
                5220: data_o = 32'h00000000 /* 0x5190 */;
                5221: data_o = 32'h00000000 /* 0x5194 */;
                5222: data_o = 32'h00000000 /* 0x5198 */;
                5223: data_o = 32'h00000000 /* 0x519c */;
                5224: data_o = 32'h00000000 /* 0x51a0 */;
                5225: data_o = 32'h00000000 /* 0x51a4 */;
                5226: data_o = 32'h00000000 /* 0x51a8 */;
                5227: data_o = 32'h00000000 /* 0x51ac */;
                5228: data_o = 32'h00000000 /* 0x51b0 */;
                5229: data_o = 32'h00000000 /* 0x51b4 */;
                5230: data_o = 32'h00000000 /* 0x51b8 */;
                5231: data_o = 32'h00000000 /* 0x51bc */;
                5232: data_o = 32'h00000000 /* 0x51c0 */;
                5233: data_o = 32'h00000000 /* 0x51c4 */;
                5234: data_o = 32'h00000000 /* 0x51c8 */;
                5235: data_o = 32'h00000000 /* 0x51cc */;
                5236: data_o = 32'h00000000 /* 0x51d0 */;
                5237: data_o = 32'h00000000 /* 0x51d4 */;
                5238: data_o = 32'h00000000 /* 0x51d8 */;
                5239: data_o = 32'h00000000 /* 0x51dc */;
                5240: data_o = 32'h00000000 /* 0x51e0 */;
                5241: data_o = 32'h00000000 /* 0x51e4 */;
                5242: data_o = 32'h00000000 /* 0x51e8 */;
                5243: data_o = 32'h00000000 /* 0x51ec */;
                5244: data_o = 32'h00000000 /* 0x51f0 */;
                5245: data_o = 32'h00000000 /* 0x51f4 */;
                5246: data_o = 32'h00000000 /* 0x51f8 */;
                5247: data_o = 32'h00000000 /* 0x51fc */;
                5248: data_o = 32'h00000000 /* 0x5200 */;
                5249: data_o = 32'h00000000 /* 0x5204 */;
                5250: data_o = 32'h00000000 /* 0x5208 */;
                5251: data_o = 32'h00000000 /* 0x520c */;
                5252: data_o = 32'h00000000 /* 0x5210 */;
                5253: data_o = 32'h00000000 /* 0x5214 */;
                5254: data_o = 32'h00000000 /* 0x5218 */;
                5255: data_o = 32'h00000000 /* 0x521c */;
                5256: data_o = 32'h00000000 /* 0x5220 */;
                5257: data_o = 32'h00000000 /* 0x5224 */;
                5258: data_o = 32'h00000000 /* 0x5228 */;
                5259: data_o = 32'h00000000 /* 0x522c */;
                5260: data_o = 32'h00000000 /* 0x5230 */;
                5261: data_o = 32'h00000000 /* 0x5234 */;
                5262: data_o = 32'h00000000 /* 0x5238 */;
                5263: data_o = 32'h00000000 /* 0x523c */;
                5264: data_o = 32'h00000000 /* 0x5240 */;
                5265: data_o = 32'h00000000 /* 0x5244 */;
                5266: data_o = 32'h00000000 /* 0x5248 */;
                5267: data_o = 32'h00000000 /* 0x524c */;
                5268: data_o = 32'h00000000 /* 0x5250 */;
                5269: data_o = 32'h00000000 /* 0x5254 */;
                5270: data_o = 32'h00000000 /* 0x5258 */;
                5271: data_o = 32'h00000000 /* 0x525c */;
                5272: data_o = 32'h00000000 /* 0x5260 */;
                5273: data_o = 32'h00000000 /* 0x5264 */;
                5274: data_o = 32'h00000000 /* 0x5268 */;
                5275: data_o = 32'h00000000 /* 0x526c */;
                5276: data_o = 32'h00000000 /* 0x5270 */;
                5277: data_o = 32'h00000000 /* 0x5274 */;
                5278: data_o = 32'h00000000 /* 0x5278 */;
                5279: data_o = 32'h00000000 /* 0x527c */;
                5280: data_o = 32'h00000000 /* 0x5280 */;
                5281: data_o = 32'h00000000 /* 0x5284 */;
                5282: data_o = 32'h00000000 /* 0x5288 */;
                5283: data_o = 32'h00000000 /* 0x528c */;
                5284: data_o = 32'h00000000 /* 0x5290 */;
                5285: data_o = 32'h00000000 /* 0x5294 */;
                5286: data_o = 32'h00000000 /* 0x5298 */;
                5287: data_o = 32'h00000000 /* 0x529c */;
                5288: data_o = 32'h00000000 /* 0x52a0 */;
                5289: data_o = 32'h00000000 /* 0x52a4 */;
                5290: data_o = 32'h00000000 /* 0x52a8 */;
                5291: data_o = 32'h00000000 /* 0x52ac */;
                5292: data_o = 32'h00000000 /* 0x52b0 */;
                5293: data_o = 32'h00000000 /* 0x52b4 */;
                5294: data_o = 32'h00000000 /* 0x52b8 */;
                5295: data_o = 32'h00000000 /* 0x52bc */;
                5296: data_o = 32'h00000000 /* 0x52c0 */;
                5297: data_o = 32'h00000000 /* 0x52c4 */;
                5298: data_o = 32'h00000000 /* 0x52c8 */;
                5299: data_o = 32'h00000000 /* 0x52cc */;
                5300: data_o = 32'h00000000 /* 0x52d0 */;
                5301: data_o = 32'h00000000 /* 0x52d4 */;
                5302: data_o = 32'h00000000 /* 0x52d8 */;
                5303: data_o = 32'h00000000 /* 0x52dc */;
                5304: data_o = 32'h00000000 /* 0x52e0 */;
                5305: data_o = 32'h00000000 /* 0x52e4 */;
                5306: data_o = 32'h00000000 /* 0x52e8 */;
                5307: data_o = 32'h00000000 /* 0x52ec */;
                5308: data_o = 32'h00000000 /* 0x52f0 */;
                5309: data_o = 32'h00000000 /* 0x52f4 */;
                5310: data_o = 32'h00000000 /* 0x52f8 */;
                5311: data_o = 32'h00000000 /* 0x52fc */;
                5312: data_o = 32'h00000000 /* 0x5300 */;
                5313: data_o = 32'h00000000 /* 0x5304 */;
                5314: data_o = 32'h00000000 /* 0x5308 */;
                5315: data_o = 32'h00000000 /* 0x530c */;
                5316: data_o = 32'h00000000 /* 0x5310 */;
                5317: data_o = 32'h00000000 /* 0x5314 */;
                5318: data_o = 32'h00000000 /* 0x5318 */;
                5319: data_o = 32'h00000000 /* 0x531c */;
                5320: data_o = 32'h00000000 /* 0x5320 */;
                5321: data_o = 32'h00000000 /* 0x5324 */;
                5322: data_o = 32'h00000000 /* 0x5328 */;
                5323: data_o = 32'h00000000 /* 0x532c */;
                5324: data_o = 32'h00000000 /* 0x5330 */;
                5325: data_o = 32'h00000000 /* 0x5334 */;
                5326: data_o = 32'h00000000 /* 0x5338 */;
                5327: data_o = 32'h00000000 /* 0x533c */;
                5328: data_o = 32'h00000000 /* 0x5340 */;
                5329: data_o = 32'h00000000 /* 0x5344 */;
                5330: data_o = 32'h00000000 /* 0x5348 */;
                5331: data_o = 32'h00000000 /* 0x534c */;
                5332: data_o = 32'h00000000 /* 0x5350 */;
                5333: data_o = 32'h00000000 /* 0x5354 */;
                5334: data_o = 32'h00000000 /* 0x5358 */;
                5335: data_o = 32'h00000000 /* 0x535c */;
                5336: data_o = 32'h00000000 /* 0x5360 */;
                5337: data_o = 32'h00000000 /* 0x5364 */;
                5338: data_o = 32'h00000000 /* 0x5368 */;
                5339: data_o = 32'h00000000 /* 0x536c */;
                5340: data_o = 32'h00000000 /* 0x5370 */;
                5341: data_o = 32'h00000000 /* 0x5374 */;
                5342: data_o = 32'h00000000 /* 0x5378 */;
                5343: data_o = 32'h00000000 /* 0x537c */;
                5344: data_o = 32'h00000000 /* 0x5380 */;
                5345: data_o = 32'h00000000 /* 0x5384 */;
                5346: data_o = 32'h00000000 /* 0x5388 */;
                5347: data_o = 32'h00000000 /* 0x538c */;
                5348: data_o = 32'h00000000 /* 0x5390 */;
                5349: data_o = 32'h00000000 /* 0x5394 */;
                5350: data_o = 32'h00000000 /* 0x5398 */;
                5351: data_o = 32'h00000000 /* 0x539c */;
                5352: data_o = 32'h00000000 /* 0x53a0 */;
                5353: data_o = 32'h00000000 /* 0x53a4 */;
                5354: data_o = 32'h00000000 /* 0x53a8 */;
                5355: data_o = 32'h00000000 /* 0x53ac */;
                5356: data_o = 32'h00000000 /* 0x53b0 */;
                5357: data_o = 32'h00000000 /* 0x53b4 */;
                5358: data_o = 32'h00000000 /* 0x53b8 */;
                5359: data_o = 32'h00000000 /* 0x53bc */;
                5360: data_o = 32'h00000000 /* 0x53c0 */;
                5361: data_o = 32'h00000000 /* 0x53c4 */;
                5362: data_o = 32'h00000000 /* 0x53c8 */;
                5363: data_o = 32'h00000000 /* 0x53cc */;
                5364: data_o = 32'h00000000 /* 0x53d0 */;
                5365: data_o = 32'h00000000 /* 0x53d4 */;
                5366: data_o = 32'h00000000 /* 0x53d8 */;
                5367: data_o = 32'h00000000 /* 0x53dc */;
                5368: data_o = 32'h00000000 /* 0x53e0 */;
                5369: data_o = 32'h00000000 /* 0x53e4 */;
                5370: data_o = 32'h00000000 /* 0x53e8 */;
                5371: data_o = 32'h00000000 /* 0x53ec */;
                5372: data_o = 32'h00000000 /* 0x53f0 */;
                5373: data_o = 32'h00000000 /* 0x53f4 */;
                5374: data_o = 32'h00000000 /* 0x53f8 */;
                5375: data_o = 32'h00000000 /* 0x53fc */;
                5376: data_o = 32'h00000000 /* 0x5400 */;
                5377: data_o = 32'h00000000 /* 0x5404 */;
                5378: data_o = 32'h00000000 /* 0x5408 */;
                5379: data_o = 32'h00000000 /* 0x540c */;
                5380: data_o = 32'h00000000 /* 0x5410 */;
                5381: data_o = 32'h00000000 /* 0x5414 */;
                5382: data_o = 32'h00000000 /* 0x5418 */;
                5383: data_o = 32'h00000000 /* 0x541c */;
                5384: data_o = 32'h00000000 /* 0x5420 */;
                5385: data_o = 32'h00000000 /* 0x5424 */;
                5386: data_o = 32'h00000000 /* 0x5428 */;
                5387: data_o = 32'h00000000 /* 0x542c */;
                5388: data_o = 32'h00000000 /* 0x5430 */;
                5389: data_o = 32'h00000000 /* 0x5434 */;
                5390: data_o = 32'h00000000 /* 0x5438 */;
                5391: data_o = 32'h00000000 /* 0x543c */;
                5392: data_o = 32'h00000000 /* 0x5440 */;
                5393: data_o = 32'h00000000 /* 0x5444 */;
                5394: data_o = 32'h00000000 /* 0x5448 */;
                5395: data_o = 32'h00000000 /* 0x544c */;
                5396: data_o = 32'h00000000 /* 0x5450 */;
                5397: data_o = 32'h00000000 /* 0x5454 */;
                5398: data_o = 32'h00000000 /* 0x5458 */;
                5399: data_o = 32'h00000000 /* 0x545c */;
                5400: data_o = 32'h00000000 /* 0x5460 */;
                5401: data_o = 32'h00000000 /* 0x5464 */;
                5402: data_o = 32'h00000000 /* 0x5468 */;
                5403: data_o = 32'h00000000 /* 0x546c */;
                5404: data_o = 32'h00000000 /* 0x5470 */;
                5405: data_o = 32'h00000000 /* 0x5474 */;
                5406: data_o = 32'h00000000 /* 0x5478 */;
                5407: data_o = 32'h00000000 /* 0x547c */;
                5408: data_o = 32'h00000000 /* 0x5480 */;
                5409: data_o = 32'h00000000 /* 0x5484 */;
                5410: data_o = 32'h00000000 /* 0x5488 */;
                5411: data_o = 32'h00000000 /* 0x548c */;
                5412: data_o = 32'h00000000 /* 0x5490 */;
                5413: data_o = 32'h00000000 /* 0x5494 */;
                5414: data_o = 32'h00000000 /* 0x5498 */;
                5415: data_o = 32'h00000000 /* 0x549c */;
                5416: data_o = 32'h00000000 /* 0x54a0 */;
                5417: data_o = 32'h00000000 /* 0x54a4 */;
                5418: data_o = 32'h00000000 /* 0x54a8 */;
                5419: data_o = 32'h00000000 /* 0x54ac */;
                5420: data_o = 32'h00000000 /* 0x54b0 */;
                5421: data_o = 32'h00000000 /* 0x54b4 */;
                5422: data_o = 32'h00000000 /* 0x54b8 */;
                5423: data_o = 32'h00000000 /* 0x54bc */;
                5424: data_o = 32'h00000000 /* 0x54c0 */;
                5425: data_o = 32'h00000000 /* 0x54c4 */;
                5426: data_o = 32'h00000000 /* 0x54c8 */;
                5427: data_o = 32'h00000000 /* 0x54cc */;
                5428: data_o = 32'h00000000 /* 0x54d0 */;
                5429: data_o = 32'h00000000 /* 0x54d4 */;
                5430: data_o = 32'h00000000 /* 0x54d8 */;
                5431: data_o = 32'h00000000 /* 0x54dc */;
                5432: data_o = 32'h00000000 /* 0x54e0 */;
                5433: data_o = 32'h00000000 /* 0x54e4 */;
                5434: data_o = 32'h00000000 /* 0x54e8 */;
                5435: data_o = 32'h00000000 /* 0x54ec */;
                5436: data_o = 32'h00000000 /* 0x54f0 */;
                5437: data_o = 32'h00000000 /* 0x54f4 */;
                5438: data_o = 32'h00000000 /* 0x54f8 */;
                5439: data_o = 32'h00000000 /* 0x54fc */;
                5440: data_o = 32'h00000000 /* 0x5500 */;
                5441: data_o = 32'h00000000 /* 0x5504 */;
                5442: data_o = 32'h00000000 /* 0x5508 */;
                5443: data_o = 32'h00000000 /* 0x550c */;
                5444: data_o = 32'h00000000 /* 0x5510 */;
                5445: data_o = 32'h00000000 /* 0x5514 */;
                5446: data_o = 32'h00000000 /* 0x5518 */;
                5447: data_o = 32'h00000000 /* 0x551c */;
                5448: data_o = 32'h00000000 /* 0x5520 */;
                5449: data_o = 32'h00000000 /* 0x5524 */;
                5450: data_o = 32'h00000000 /* 0x5528 */;
                5451: data_o = 32'h00000000 /* 0x552c */;
                5452: data_o = 32'h00000000 /* 0x5530 */;
                5453: data_o = 32'h00000000 /* 0x5534 */;
                5454: data_o = 32'h00000000 /* 0x5538 */;
                5455: data_o = 32'h00000000 /* 0x553c */;
                5456: data_o = 32'h00000000 /* 0x5540 */;
                5457: data_o = 32'h00000000 /* 0x5544 */;
                5458: data_o = 32'h00000000 /* 0x5548 */;
                5459: data_o = 32'h00000000 /* 0x554c */;
                5460: data_o = 32'h00000000 /* 0x5550 */;
                5461: data_o = 32'h00000000 /* 0x5554 */;
                5462: data_o = 32'h00000000 /* 0x5558 */;
                5463: data_o = 32'h00000000 /* 0x555c */;
                5464: data_o = 32'h00000000 /* 0x5560 */;
                5465: data_o = 32'h00000000 /* 0x5564 */;
                5466: data_o = 32'h00000000 /* 0x5568 */;
                5467: data_o = 32'h00000000 /* 0x556c */;
                5468: data_o = 32'h00000000 /* 0x5570 */;
                5469: data_o = 32'h00000000 /* 0x5574 */;
                5470: data_o = 32'h00000000 /* 0x5578 */;
                5471: data_o = 32'h00000000 /* 0x557c */;
                5472: data_o = 32'h00000000 /* 0x5580 */;
                5473: data_o = 32'h00000000 /* 0x5584 */;
                5474: data_o = 32'h00000000 /* 0x5588 */;
                5475: data_o = 32'h00000000 /* 0x558c */;
                5476: data_o = 32'h00000000 /* 0x5590 */;
                5477: data_o = 32'h00000000 /* 0x5594 */;
                5478: data_o = 32'h00000000 /* 0x5598 */;
                5479: data_o = 32'h00000000 /* 0x559c */;
                5480: data_o = 32'h00000000 /* 0x55a0 */;
                5481: data_o = 32'h00000000 /* 0x55a4 */;
                5482: data_o = 32'h00000000 /* 0x55a8 */;
                5483: data_o = 32'h00000000 /* 0x55ac */;
                5484: data_o = 32'h00000000 /* 0x55b0 */;
                5485: data_o = 32'h00000000 /* 0x55b4 */;
                5486: data_o = 32'h00000000 /* 0x55b8 */;
                5487: data_o = 32'h00000000 /* 0x55bc */;
                5488: data_o = 32'h00000000 /* 0x55c0 */;
                5489: data_o = 32'h00000000 /* 0x55c4 */;
                5490: data_o = 32'h00000000 /* 0x55c8 */;
                5491: data_o = 32'h00000000 /* 0x55cc */;
                5492: data_o = 32'h00000000 /* 0x55d0 */;
                5493: data_o = 32'h00000000 /* 0x55d4 */;
                5494: data_o = 32'h00000000 /* 0x55d8 */;
                5495: data_o = 32'h00000000 /* 0x55dc */;
                5496: data_o = 32'h00000000 /* 0x55e0 */;
                5497: data_o = 32'h00000000 /* 0x55e4 */;
                5498: data_o = 32'h00000000 /* 0x55e8 */;
                5499: data_o = 32'h00000000 /* 0x55ec */;
                5500: data_o = 32'h00000000 /* 0x55f0 */;
                5501: data_o = 32'h00000000 /* 0x55f4 */;
                5502: data_o = 32'h00000000 /* 0x55f8 */;
                5503: data_o = 32'h00000000 /* 0x55fc */;
                5504: data_o = 32'h00000000 /* 0x5600 */;
                5505: data_o = 32'h00000000 /* 0x5604 */;
                5506: data_o = 32'h00000000 /* 0x5608 */;
                5507: data_o = 32'h00000000 /* 0x560c */;
                5508: data_o = 32'h00000000 /* 0x5610 */;
                5509: data_o = 32'h00000000 /* 0x5614 */;
                5510: data_o = 32'h00000000 /* 0x5618 */;
                5511: data_o = 32'h00000000 /* 0x561c */;
                5512: data_o = 32'h00000000 /* 0x5620 */;
                5513: data_o = 32'h00000000 /* 0x5624 */;
                5514: data_o = 32'h00000000 /* 0x5628 */;
                5515: data_o = 32'h00000000 /* 0x562c */;
                5516: data_o = 32'h00000000 /* 0x5630 */;
                5517: data_o = 32'h00000000 /* 0x5634 */;
                5518: data_o = 32'h00000000 /* 0x5638 */;
                5519: data_o = 32'h00000000 /* 0x563c */;
                5520: data_o = 32'h00000000 /* 0x5640 */;
                5521: data_o = 32'h00000000 /* 0x5644 */;
                5522: data_o = 32'h00000000 /* 0x5648 */;
                5523: data_o = 32'h00000000 /* 0x564c */;
                5524: data_o = 32'h00000000 /* 0x5650 */;
                5525: data_o = 32'h00000000 /* 0x5654 */;
                5526: data_o = 32'h00000000 /* 0x5658 */;
                5527: data_o = 32'h00000000 /* 0x565c */;
                5528: data_o = 32'h00000000 /* 0x5660 */;
                5529: data_o = 32'h00000000 /* 0x5664 */;
                5530: data_o = 32'h00000000 /* 0x5668 */;
                5531: data_o = 32'h00000000 /* 0x566c */;
                5532: data_o = 32'h00000000 /* 0x5670 */;
                5533: data_o = 32'h00000000 /* 0x5674 */;
                5534: data_o = 32'h00000000 /* 0x5678 */;
                5535: data_o = 32'h00000000 /* 0x567c */;
                5536: data_o = 32'h00000000 /* 0x5680 */;
                5537: data_o = 32'h00000000 /* 0x5684 */;
                5538: data_o = 32'h00000000 /* 0x5688 */;
                5539: data_o = 32'h00000000 /* 0x568c */;
                5540: data_o = 32'h00000000 /* 0x5690 */;
                5541: data_o = 32'h00000000 /* 0x5694 */;
                5542: data_o = 32'h00000000 /* 0x5698 */;
                5543: data_o = 32'h00000000 /* 0x569c */;
                5544: data_o = 32'h00000000 /* 0x56a0 */;
                5545: data_o = 32'h00000000 /* 0x56a4 */;
                5546: data_o = 32'h00000000 /* 0x56a8 */;
                5547: data_o = 32'h00000000 /* 0x56ac */;
                5548: data_o = 32'h00000000 /* 0x56b0 */;
                5549: data_o = 32'h00000000 /* 0x56b4 */;
                5550: data_o = 32'h00000000 /* 0x56b8 */;
                5551: data_o = 32'h00000000 /* 0x56bc */;
                5552: data_o = 32'h00000000 /* 0x56c0 */;
                5553: data_o = 32'h00000000 /* 0x56c4 */;
                5554: data_o = 32'h00000000 /* 0x56c8 */;
                5555: data_o = 32'h00000000 /* 0x56cc */;
                5556: data_o = 32'h00000000 /* 0x56d0 */;
                5557: data_o = 32'h00000000 /* 0x56d4 */;
                5558: data_o = 32'h00000000 /* 0x56d8 */;
                5559: data_o = 32'h00000000 /* 0x56dc */;
                5560: data_o = 32'h00000000 /* 0x56e0 */;
                5561: data_o = 32'h00000000 /* 0x56e4 */;
                5562: data_o = 32'h00000000 /* 0x56e8 */;
                5563: data_o = 32'h00000000 /* 0x56ec */;
                5564: data_o = 32'h00000000 /* 0x56f0 */;
                5565: data_o = 32'h00000000 /* 0x56f4 */;
                5566: data_o = 32'h00000000 /* 0x56f8 */;
                5567: data_o = 32'h00000000 /* 0x56fc */;
                5568: data_o = 32'h00000000 /* 0x5700 */;
                5569: data_o = 32'h00000000 /* 0x5704 */;
                5570: data_o = 32'h00000000 /* 0x5708 */;
                5571: data_o = 32'h00000000 /* 0x570c */;
                5572: data_o = 32'h00000000 /* 0x5710 */;
                5573: data_o = 32'h00000000 /* 0x5714 */;
                5574: data_o = 32'h00000000 /* 0x5718 */;
                5575: data_o = 32'h00000000 /* 0x571c */;
                5576: data_o = 32'h00000000 /* 0x5720 */;
                5577: data_o = 32'h00000000 /* 0x5724 */;
                5578: data_o = 32'h00000000 /* 0x5728 */;
                5579: data_o = 32'h00000000 /* 0x572c */;
                5580: data_o = 32'h00000000 /* 0x5730 */;
                5581: data_o = 32'h00000000 /* 0x5734 */;
                5582: data_o = 32'h00000000 /* 0x5738 */;
                5583: data_o = 32'h00000000 /* 0x573c */;
                5584: data_o = 32'h00000000 /* 0x5740 */;
                5585: data_o = 32'h00000000 /* 0x5744 */;
                5586: data_o = 32'h00000000 /* 0x5748 */;
                5587: data_o = 32'h00000000 /* 0x574c */;
                5588: data_o = 32'h00000000 /* 0x5750 */;
                5589: data_o = 32'h00000000 /* 0x5754 */;
                5590: data_o = 32'h00000000 /* 0x5758 */;
                5591: data_o = 32'h00000000 /* 0x575c */;
                5592: data_o = 32'h00000000 /* 0x5760 */;
                5593: data_o = 32'h00000000 /* 0x5764 */;
                5594: data_o = 32'h00000000 /* 0x5768 */;
                5595: data_o = 32'h00000000 /* 0x576c */;
                5596: data_o = 32'h00000000 /* 0x5770 */;
                5597: data_o = 32'h00000000 /* 0x5774 */;
                5598: data_o = 32'h00000000 /* 0x5778 */;
                5599: data_o = 32'h00000000 /* 0x577c */;
                5600: data_o = 32'h00000000 /* 0x5780 */;
                5601: data_o = 32'h00000000 /* 0x5784 */;
                5602: data_o = 32'h00000000 /* 0x5788 */;
                5603: data_o = 32'h00000000 /* 0x578c */;
                5604: data_o = 32'h00000000 /* 0x5790 */;
                5605: data_o = 32'h00000000 /* 0x5794 */;
                5606: data_o = 32'h00000000 /* 0x5798 */;
                5607: data_o = 32'h00000000 /* 0x579c */;
                5608: data_o = 32'h00000000 /* 0x57a0 */;
                5609: data_o = 32'h00000000 /* 0x57a4 */;
                5610: data_o = 32'h00000000 /* 0x57a8 */;
                5611: data_o = 32'h00000000 /* 0x57ac */;
                5612: data_o = 32'h00000000 /* 0x57b0 */;
                5613: data_o = 32'h00000000 /* 0x57b4 */;
                5614: data_o = 32'h00000000 /* 0x57b8 */;
                5615: data_o = 32'h00000000 /* 0x57bc */;
                5616: data_o = 32'h00000000 /* 0x57c0 */;
                5617: data_o = 32'h00000000 /* 0x57c4 */;
                5618: data_o = 32'h00000000 /* 0x57c8 */;
                5619: data_o = 32'h00000000 /* 0x57cc */;
                5620: data_o = 32'h00000000 /* 0x57d0 */;
                5621: data_o = 32'h00000000 /* 0x57d4 */;
                5622: data_o = 32'h00000000 /* 0x57d8 */;
                5623: data_o = 32'h00000000 /* 0x57dc */;
                5624: data_o = 32'h00000000 /* 0x57e0 */;
                5625: data_o = 32'h00000000 /* 0x57e4 */;
                5626: data_o = 32'h00000000 /* 0x57e8 */;
                5627: data_o = 32'h00000000 /* 0x57ec */;
                5628: data_o = 32'h00000000 /* 0x57f0 */;
                5629: data_o = 32'h00000000 /* 0x57f4 */;
                5630: data_o = 32'h00000000 /* 0x57f8 */;
                5631: data_o = 32'h00000000 /* 0x57fc */;
                5632: data_o = 32'h00000000 /* 0x5800 */;
                5633: data_o = 32'h00000000 /* 0x5804 */;
                5634: data_o = 32'h00000000 /* 0x5808 */;
                5635: data_o = 32'h00000000 /* 0x580c */;
                5636: data_o = 32'h00000000 /* 0x5810 */;
                5637: data_o = 32'h00000000 /* 0x5814 */;
                5638: data_o = 32'h00000000 /* 0x5818 */;
                5639: data_o = 32'h00000000 /* 0x581c */;
                5640: data_o = 32'h00000000 /* 0x5820 */;
                5641: data_o = 32'h00000000 /* 0x5824 */;
                5642: data_o = 32'h00000000 /* 0x5828 */;
                5643: data_o = 32'h00000000 /* 0x582c */;
                5644: data_o = 32'h00000000 /* 0x5830 */;
                5645: data_o = 32'h00000000 /* 0x5834 */;
                5646: data_o = 32'h00000000 /* 0x5838 */;
                5647: data_o = 32'h00000000 /* 0x583c */;
                5648: data_o = 32'h00000000 /* 0x5840 */;
                5649: data_o = 32'h00000000 /* 0x5844 */;
                5650: data_o = 32'h00000000 /* 0x5848 */;
                5651: data_o = 32'h00000000 /* 0x584c */;
                5652: data_o = 32'h00000000 /* 0x5850 */;
                5653: data_o = 32'h00000000 /* 0x5854 */;
                5654: data_o = 32'h00000000 /* 0x5858 */;
                5655: data_o = 32'h00000000 /* 0x585c */;
                5656: data_o = 32'h00000000 /* 0x5860 */;
                5657: data_o = 32'h00000000 /* 0x5864 */;
                5658: data_o = 32'h00000000 /* 0x5868 */;
                5659: data_o = 32'h00000000 /* 0x586c */;
                5660: data_o = 32'h00000000 /* 0x5870 */;
                5661: data_o = 32'h00000000 /* 0x5874 */;
                5662: data_o = 32'h00000000 /* 0x5878 */;
                5663: data_o = 32'h00000000 /* 0x587c */;
                5664: data_o = 32'h00000000 /* 0x5880 */;
                5665: data_o = 32'h00000000 /* 0x5884 */;
                5666: data_o = 32'h00000000 /* 0x5888 */;
                5667: data_o = 32'h00000000 /* 0x588c */;
                5668: data_o = 32'h00000000 /* 0x5890 */;
                5669: data_o = 32'h00000000 /* 0x5894 */;
                5670: data_o = 32'h00000000 /* 0x5898 */;
                5671: data_o = 32'h00000000 /* 0x589c */;
                5672: data_o = 32'h00000000 /* 0x58a0 */;
                5673: data_o = 32'h00000000 /* 0x58a4 */;
                5674: data_o = 32'h00000000 /* 0x58a8 */;
                5675: data_o = 32'h00000000 /* 0x58ac */;
                5676: data_o = 32'h00000000 /* 0x58b0 */;
                5677: data_o = 32'h00000000 /* 0x58b4 */;
                5678: data_o = 32'h00000000 /* 0x58b8 */;
                5679: data_o = 32'h00000000 /* 0x58bc */;
                5680: data_o = 32'h00000000 /* 0x58c0 */;
                5681: data_o = 32'h00000000 /* 0x58c4 */;
                5682: data_o = 32'h00000000 /* 0x58c8 */;
                5683: data_o = 32'h00000000 /* 0x58cc */;
                5684: data_o = 32'h00000000 /* 0x58d0 */;
                5685: data_o = 32'h00000000 /* 0x58d4 */;
                5686: data_o = 32'h00000000 /* 0x58d8 */;
                5687: data_o = 32'h00000000 /* 0x58dc */;
                5688: data_o = 32'h00000000 /* 0x58e0 */;
                5689: data_o = 32'h00000000 /* 0x58e4 */;
                5690: data_o = 32'h00000000 /* 0x58e8 */;
                5691: data_o = 32'h00000000 /* 0x58ec */;
                5692: data_o = 32'h00000000 /* 0x58f0 */;
                5693: data_o = 32'h00000000 /* 0x58f4 */;
                5694: data_o = 32'h00000000 /* 0x58f8 */;
                5695: data_o = 32'h00000000 /* 0x58fc */;
                5696: data_o = 32'h00000000 /* 0x5900 */;
                5697: data_o = 32'h00000000 /* 0x5904 */;
                5698: data_o = 32'h00000000 /* 0x5908 */;
                5699: data_o = 32'h00000000 /* 0x590c */;
                5700: data_o = 32'h00000000 /* 0x5910 */;
                5701: data_o = 32'h00000000 /* 0x5914 */;
                5702: data_o = 32'h00000000 /* 0x5918 */;
                5703: data_o = 32'h00000000 /* 0x591c */;
                5704: data_o = 32'h00000000 /* 0x5920 */;
                5705: data_o = 32'h00000000 /* 0x5924 */;
                5706: data_o = 32'h00000000 /* 0x5928 */;
                5707: data_o = 32'h00000000 /* 0x592c */;
                5708: data_o = 32'h00000000 /* 0x5930 */;
                5709: data_o = 32'h00000000 /* 0x5934 */;
                5710: data_o = 32'h00000000 /* 0x5938 */;
                5711: data_o = 32'h00000000 /* 0x593c */;
                5712: data_o = 32'h00000000 /* 0x5940 */;
                5713: data_o = 32'h00000000 /* 0x5944 */;
                5714: data_o = 32'h00000000 /* 0x5948 */;
                5715: data_o = 32'h00000000 /* 0x594c */;
                5716: data_o = 32'h00000000 /* 0x5950 */;
                5717: data_o = 32'h00000000 /* 0x5954 */;
                5718: data_o = 32'h00000000 /* 0x5958 */;
                5719: data_o = 32'h00000000 /* 0x595c */;
                5720: data_o = 32'h00000000 /* 0x5960 */;
                5721: data_o = 32'h00000000 /* 0x5964 */;
                5722: data_o = 32'h00000000 /* 0x5968 */;
                5723: data_o = 32'h00000000 /* 0x596c */;
                5724: data_o = 32'h00000000 /* 0x5970 */;
                5725: data_o = 32'h00000000 /* 0x5974 */;
                5726: data_o = 32'h00000000 /* 0x5978 */;
                5727: data_o = 32'h00000000 /* 0x597c */;
                5728: data_o = 32'h00000000 /* 0x5980 */;
                5729: data_o = 32'h00000000 /* 0x5984 */;
                5730: data_o = 32'h00000000 /* 0x5988 */;
                5731: data_o = 32'h00000000 /* 0x598c */;
                5732: data_o = 32'h00000000 /* 0x5990 */;
                5733: data_o = 32'h00000000 /* 0x5994 */;
                5734: data_o = 32'h00000000 /* 0x5998 */;
                5735: data_o = 32'h00000000 /* 0x599c */;
                5736: data_o = 32'h00000000 /* 0x59a0 */;
                5737: data_o = 32'h00000000 /* 0x59a4 */;
                5738: data_o = 32'h00000000 /* 0x59a8 */;
                5739: data_o = 32'h00000000 /* 0x59ac */;
                5740: data_o = 32'h00000000 /* 0x59b0 */;
                5741: data_o = 32'h00000000 /* 0x59b4 */;
                5742: data_o = 32'h00000000 /* 0x59b8 */;
                5743: data_o = 32'h00000000 /* 0x59bc */;
                5744: data_o = 32'h00000000 /* 0x59c0 */;
                5745: data_o = 32'h00000000 /* 0x59c4 */;
                5746: data_o = 32'h00000000 /* 0x59c8 */;
                5747: data_o = 32'h00000000 /* 0x59cc */;
                5748: data_o = 32'h00000000 /* 0x59d0 */;
                5749: data_o = 32'h00000000 /* 0x59d4 */;
                5750: data_o = 32'h00000000 /* 0x59d8 */;
                5751: data_o = 32'h00000000 /* 0x59dc */;
                5752: data_o = 32'h00000000 /* 0x59e0 */;
                5753: data_o = 32'h00000000 /* 0x59e4 */;
                5754: data_o = 32'h00000000 /* 0x59e8 */;
                5755: data_o = 32'h00000000 /* 0x59ec */;
                5756: data_o = 32'h00000000 /* 0x59f0 */;
                5757: data_o = 32'h00000000 /* 0x59f4 */;
                5758: data_o = 32'h00000000 /* 0x59f8 */;
                5759: data_o = 32'h00000000 /* 0x59fc */;
                5760: data_o = 32'h00000000 /* 0x5a00 */;
                5761: data_o = 32'h00000000 /* 0x5a04 */;
                5762: data_o = 32'h00000000 /* 0x5a08 */;
                5763: data_o = 32'h00000000 /* 0x5a0c */;
                5764: data_o = 32'h00000000 /* 0x5a10 */;
                5765: data_o = 32'h00000000 /* 0x5a14 */;
                5766: data_o = 32'h00000000 /* 0x5a18 */;
                5767: data_o = 32'h00000000 /* 0x5a1c */;
                5768: data_o = 32'h00000000 /* 0x5a20 */;
                5769: data_o = 32'h00000000 /* 0x5a24 */;
                5770: data_o = 32'h00000000 /* 0x5a28 */;
                5771: data_o = 32'h00000000 /* 0x5a2c */;
                5772: data_o = 32'h00000000 /* 0x5a30 */;
                5773: data_o = 32'h00000000 /* 0x5a34 */;
                5774: data_o = 32'h00000000 /* 0x5a38 */;
                5775: data_o = 32'h00000000 /* 0x5a3c */;
                5776: data_o = 32'h00000000 /* 0x5a40 */;
                5777: data_o = 32'h00000000 /* 0x5a44 */;
                5778: data_o = 32'h00000000 /* 0x5a48 */;
                5779: data_o = 32'h00000000 /* 0x5a4c */;
                5780: data_o = 32'h00000000 /* 0x5a50 */;
                5781: data_o = 32'h00000000 /* 0x5a54 */;
                5782: data_o = 32'h00000000 /* 0x5a58 */;
                5783: data_o = 32'h00000000 /* 0x5a5c */;
                5784: data_o = 32'h00000000 /* 0x5a60 */;
                5785: data_o = 32'h00000000 /* 0x5a64 */;
                5786: data_o = 32'h00000000 /* 0x5a68 */;
                5787: data_o = 32'h00000000 /* 0x5a6c */;
                5788: data_o = 32'h00000000 /* 0x5a70 */;
                5789: data_o = 32'h00000000 /* 0x5a74 */;
                5790: data_o = 32'h00000000 /* 0x5a78 */;
                5791: data_o = 32'h00000000 /* 0x5a7c */;
                5792: data_o = 32'h00000000 /* 0x5a80 */;
                5793: data_o = 32'h00000000 /* 0x5a84 */;
                5794: data_o = 32'h00000000 /* 0x5a88 */;
                5795: data_o = 32'h00000000 /* 0x5a8c */;
                5796: data_o = 32'h00000000 /* 0x5a90 */;
                5797: data_o = 32'h00000000 /* 0x5a94 */;
                5798: data_o = 32'h00000000 /* 0x5a98 */;
                5799: data_o = 32'h00000000 /* 0x5a9c */;
                5800: data_o = 32'h00000000 /* 0x5aa0 */;
                5801: data_o = 32'h00000000 /* 0x5aa4 */;
                5802: data_o = 32'h00000000 /* 0x5aa8 */;
                5803: data_o = 32'h00000000 /* 0x5aac */;
                5804: data_o = 32'h00000000 /* 0x5ab0 */;
                5805: data_o = 32'h00000000 /* 0x5ab4 */;
                5806: data_o = 32'h00000000 /* 0x5ab8 */;
                5807: data_o = 32'h00000000 /* 0x5abc */;
                5808: data_o = 32'h00000000 /* 0x5ac0 */;
                5809: data_o = 32'h00000000 /* 0x5ac4 */;
                5810: data_o = 32'h00000000 /* 0x5ac8 */;
                5811: data_o = 32'h00000000 /* 0x5acc */;
                5812: data_o = 32'h00000000 /* 0x5ad0 */;
                5813: data_o = 32'h00000000 /* 0x5ad4 */;
                5814: data_o = 32'h00000000 /* 0x5ad8 */;
                5815: data_o = 32'h00000000 /* 0x5adc */;
                5816: data_o = 32'h00000000 /* 0x5ae0 */;
                5817: data_o = 32'h00000000 /* 0x5ae4 */;
                5818: data_o = 32'h00000000 /* 0x5ae8 */;
                5819: data_o = 32'h00000000 /* 0x5aec */;
                5820: data_o = 32'h00000000 /* 0x5af0 */;
                5821: data_o = 32'h00000000 /* 0x5af4 */;
                5822: data_o = 32'h00000000 /* 0x5af8 */;
                5823: data_o = 32'h00000000 /* 0x5afc */;
                5824: data_o = 32'h00000000 /* 0x5b00 */;
                5825: data_o = 32'h00000000 /* 0x5b04 */;
                5826: data_o = 32'h00000000 /* 0x5b08 */;
                5827: data_o = 32'h00000000 /* 0x5b0c */;
                5828: data_o = 32'h00000000 /* 0x5b10 */;
                5829: data_o = 32'h00000000 /* 0x5b14 */;
                5830: data_o = 32'h00000000 /* 0x5b18 */;
                5831: data_o = 32'h00000000 /* 0x5b1c */;
                5832: data_o = 32'h00000000 /* 0x5b20 */;
                5833: data_o = 32'h00000000 /* 0x5b24 */;
                5834: data_o = 32'h00000000 /* 0x5b28 */;
                5835: data_o = 32'h00000000 /* 0x5b2c */;
                5836: data_o = 32'h00000000 /* 0x5b30 */;
                5837: data_o = 32'h00000000 /* 0x5b34 */;
                5838: data_o = 32'h00000000 /* 0x5b38 */;
                5839: data_o = 32'h00000000 /* 0x5b3c */;
                5840: data_o = 32'h00000000 /* 0x5b40 */;
                5841: data_o = 32'h00000000 /* 0x5b44 */;
                5842: data_o = 32'h00000000 /* 0x5b48 */;
                5843: data_o = 32'h00000000 /* 0x5b4c */;
                5844: data_o = 32'h00000000 /* 0x5b50 */;
                5845: data_o = 32'h00000000 /* 0x5b54 */;
                5846: data_o = 32'h00000000 /* 0x5b58 */;
                5847: data_o = 32'h00000000 /* 0x5b5c */;
                5848: data_o = 32'h00000000 /* 0x5b60 */;
                5849: data_o = 32'h00000000 /* 0x5b64 */;
                5850: data_o = 32'h00000000 /* 0x5b68 */;
                5851: data_o = 32'h00000000 /* 0x5b6c */;
                5852: data_o = 32'h00000000 /* 0x5b70 */;
                5853: data_o = 32'h00000000 /* 0x5b74 */;
                5854: data_o = 32'h00000000 /* 0x5b78 */;
                5855: data_o = 32'h00000000 /* 0x5b7c */;
                5856: data_o = 32'h00000000 /* 0x5b80 */;
                5857: data_o = 32'h00000000 /* 0x5b84 */;
                5858: data_o = 32'h00000000 /* 0x5b88 */;
                5859: data_o = 32'h00000000 /* 0x5b8c */;
                5860: data_o = 32'h00000000 /* 0x5b90 */;
                5861: data_o = 32'h00000000 /* 0x5b94 */;
                5862: data_o = 32'h00000000 /* 0x5b98 */;
                5863: data_o = 32'h00000000 /* 0x5b9c */;
                5864: data_o = 32'h00000000 /* 0x5ba0 */;
                5865: data_o = 32'h00000000 /* 0x5ba4 */;
                5866: data_o = 32'h00000000 /* 0x5ba8 */;
                5867: data_o = 32'h00000000 /* 0x5bac */;
                5868: data_o = 32'h00000000 /* 0x5bb0 */;
                5869: data_o = 32'h00000000 /* 0x5bb4 */;
                5870: data_o = 32'h00000000 /* 0x5bb8 */;
                5871: data_o = 32'h00000000 /* 0x5bbc */;
                5872: data_o = 32'h00000000 /* 0x5bc0 */;
                5873: data_o = 32'h00000000 /* 0x5bc4 */;
                5874: data_o = 32'h00000000 /* 0x5bc8 */;
                5875: data_o = 32'h00000000 /* 0x5bcc */;
                5876: data_o = 32'h00000000 /* 0x5bd0 */;
                5877: data_o = 32'h00000000 /* 0x5bd4 */;
                5878: data_o = 32'h00000000 /* 0x5bd8 */;
                5879: data_o = 32'h00000000 /* 0x5bdc */;
                5880: data_o = 32'h00000000 /* 0x5be0 */;
                5881: data_o = 32'h00000000 /* 0x5be4 */;
                5882: data_o = 32'h00000000 /* 0x5be8 */;
                5883: data_o = 32'h00000000 /* 0x5bec */;
                5884: data_o = 32'h00000000 /* 0x5bf0 */;
                5885: data_o = 32'h00000000 /* 0x5bf4 */;
                5886: data_o = 32'h00000000 /* 0x5bf8 */;
                5887: data_o = 32'h00000000 /* 0x5bfc */;
                5888: data_o = 32'h00000000 /* 0x5c00 */;
                5889: data_o = 32'h00000000 /* 0x5c04 */;
                5890: data_o = 32'h00000000 /* 0x5c08 */;
                5891: data_o = 32'h00000000 /* 0x5c0c */;
                5892: data_o = 32'h00000000 /* 0x5c10 */;
                5893: data_o = 32'h00000000 /* 0x5c14 */;
                5894: data_o = 32'h00000000 /* 0x5c18 */;
                5895: data_o = 32'h00000000 /* 0x5c1c */;
                5896: data_o = 32'h00000000 /* 0x5c20 */;
                5897: data_o = 32'h00000000 /* 0x5c24 */;
                5898: data_o = 32'h00000000 /* 0x5c28 */;
                5899: data_o = 32'h00000000 /* 0x5c2c */;
                5900: data_o = 32'h00000000 /* 0x5c30 */;
                5901: data_o = 32'h00000000 /* 0x5c34 */;
                5902: data_o = 32'h00000000 /* 0x5c38 */;
                5903: data_o = 32'h00000000 /* 0x5c3c */;
                5904: data_o = 32'h00000000 /* 0x5c40 */;
                5905: data_o = 32'h00000000 /* 0x5c44 */;
                5906: data_o = 32'h00000000 /* 0x5c48 */;
                5907: data_o = 32'h00000000 /* 0x5c4c */;
                5908: data_o = 32'h00000000 /* 0x5c50 */;
                5909: data_o = 32'h00000000 /* 0x5c54 */;
                5910: data_o = 32'h00000000 /* 0x5c58 */;
                5911: data_o = 32'h00000000 /* 0x5c5c */;
                5912: data_o = 32'h00000000 /* 0x5c60 */;
                5913: data_o = 32'h00000000 /* 0x5c64 */;
                5914: data_o = 32'h00000000 /* 0x5c68 */;
                5915: data_o = 32'h00000000 /* 0x5c6c */;
                5916: data_o = 32'h00000000 /* 0x5c70 */;
                5917: data_o = 32'h00000000 /* 0x5c74 */;
                5918: data_o = 32'h00000000 /* 0x5c78 */;
                5919: data_o = 32'h00000000 /* 0x5c7c */;
                5920: data_o = 32'h00000000 /* 0x5c80 */;
                5921: data_o = 32'h00000000 /* 0x5c84 */;
                5922: data_o = 32'h00000000 /* 0x5c88 */;
                5923: data_o = 32'h00000000 /* 0x5c8c */;
                5924: data_o = 32'h00000000 /* 0x5c90 */;
                5925: data_o = 32'h00000000 /* 0x5c94 */;
                5926: data_o = 32'h00000000 /* 0x5c98 */;
                5927: data_o = 32'h00000000 /* 0x5c9c */;
                5928: data_o = 32'h00000000 /* 0x5ca0 */;
                5929: data_o = 32'h00000000 /* 0x5ca4 */;
                5930: data_o = 32'h00000000 /* 0x5ca8 */;
                5931: data_o = 32'h00000000 /* 0x5cac */;
                5932: data_o = 32'h00000000 /* 0x5cb0 */;
                5933: data_o = 32'h00000000 /* 0x5cb4 */;
                5934: data_o = 32'h00000000 /* 0x5cb8 */;
                5935: data_o = 32'h00000000 /* 0x5cbc */;
                5936: data_o = 32'h00000000 /* 0x5cc0 */;
                5937: data_o = 32'h00000000 /* 0x5cc4 */;
                5938: data_o = 32'h00000000 /* 0x5cc8 */;
                5939: data_o = 32'h00000000 /* 0x5ccc */;
                5940: data_o = 32'h00000000 /* 0x5cd0 */;
                5941: data_o = 32'h00000000 /* 0x5cd4 */;
                5942: data_o = 32'h00000000 /* 0x5cd8 */;
                5943: data_o = 32'h00000000 /* 0x5cdc */;
                5944: data_o = 32'h00000000 /* 0x5ce0 */;
                5945: data_o = 32'h00000000 /* 0x5ce4 */;
                5946: data_o = 32'h00000000 /* 0x5ce8 */;
                5947: data_o = 32'h00000000 /* 0x5cec */;
                5948: data_o = 32'h00000000 /* 0x5cf0 */;
                5949: data_o = 32'h00000000 /* 0x5cf4 */;
                5950: data_o = 32'h00000000 /* 0x5cf8 */;
                5951: data_o = 32'h00000000 /* 0x5cfc */;
                5952: data_o = 32'h00000000 /* 0x5d00 */;
                5953: data_o = 32'h00000000 /* 0x5d04 */;
                5954: data_o = 32'h00000000 /* 0x5d08 */;
                5955: data_o = 32'h00000000 /* 0x5d0c */;
                5956: data_o = 32'h00000000 /* 0x5d10 */;
                5957: data_o = 32'h00000000 /* 0x5d14 */;
                5958: data_o = 32'h00000000 /* 0x5d18 */;
                5959: data_o = 32'h00000000 /* 0x5d1c */;
                5960: data_o = 32'h00000000 /* 0x5d20 */;
                5961: data_o = 32'h00000000 /* 0x5d24 */;
                5962: data_o = 32'h00000000 /* 0x5d28 */;
                5963: data_o = 32'h00000000 /* 0x5d2c */;
                5964: data_o = 32'h00000000 /* 0x5d30 */;
                5965: data_o = 32'h00000000 /* 0x5d34 */;
                5966: data_o = 32'h00000000 /* 0x5d38 */;
                5967: data_o = 32'h00000000 /* 0x5d3c */;
                5968: data_o = 32'h00000000 /* 0x5d40 */;
                5969: data_o = 32'h00000000 /* 0x5d44 */;
                5970: data_o = 32'h00000000 /* 0x5d48 */;
                5971: data_o = 32'h00000000 /* 0x5d4c */;
                5972: data_o = 32'h00000000 /* 0x5d50 */;
                5973: data_o = 32'h00000000 /* 0x5d54 */;
                5974: data_o = 32'h00000000 /* 0x5d58 */;
                5975: data_o = 32'h00000000 /* 0x5d5c */;
                5976: data_o = 32'h00000000 /* 0x5d60 */;
                5977: data_o = 32'h00000000 /* 0x5d64 */;
                5978: data_o = 32'h00000000 /* 0x5d68 */;
                5979: data_o = 32'h00000000 /* 0x5d6c */;
                5980: data_o = 32'h00000000 /* 0x5d70 */;
                5981: data_o = 32'h00000000 /* 0x5d74 */;
                5982: data_o = 32'h00000000 /* 0x5d78 */;
                5983: data_o = 32'h00000000 /* 0x5d7c */;
                5984: data_o = 32'h00000000 /* 0x5d80 */;
                5985: data_o = 32'h00000000 /* 0x5d84 */;
                5986: data_o = 32'h00000000 /* 0x5d88 */;
                5987: data_o = 32'h00000000 /* 0x5d8c */;
                5988: data_o = 32'h00000000 /* 0x5d90 */;
                5989: data_o = 32'h00000000 /* 0x5d94 */;
                5990: data_o = 32'h00000000 /* 0x5d98 */;
                5991: data_o = 32'h00000000 /* 0x5d9c */;
                5992: data_o = 32'h00000000 /* 0x5da0 */;
                5993: data_o = 32'h00000000 /* 0x5da4 */;
                5994: data_o = 32'h00000000 /* 0x5da8 */;
                5995: data_o = 32'h00000000 /* 0x5dac */;
                5996: data_o = 32'h00000000 /* 0x5db0 */;
                5997: data_o = 32'h00000000 /* 0x5db4 */;
                5998: data_o = 32'h00000000 /* 0x5db8 */;
                5999: data_o = 32'h00000000 /* 0x5dbc */;
                6000: data_o = 32'h00000000 /* 0x5dc0 */;
                6001: data_o = 32'h00000000 /* 0x5dc4 */;
                6002: data_o = 32'h00000000 /* 0x5dc8 */;
                6003: data_o = 32'h00000000 /* 0x5dcc */;
                6004: data_o = 32'h00000000 /* 0x5dd0 */;
                6005: data_o = 32'h00000000 /* 0x5dd4 */;
                6006: data_o = 32'h00000000 /* 0x5dd8 */;
                6007: data_o = 32'h00000000 /* 0x5ddc */;
                6008: data_o = 32'h00000000 /* 0x5de0 */;
                6009: data_o = 32'h00000000 /* 0x5de4 */;
                6010: data_o = 32'h00000000 /* 0x5de8 */;
                6011: data_o = 32'h00000000 /* 0x5dec */;
                6012: data_o = 32'h00000000 /* 0x5df0 */;
                6013: data_o = 32'h00000000 /* 0x5df4 */;
                6014: data_o = 32'h00000000 /* 0x5df8 */;
                6015: data_o = 32'h00000000 /* 0x5dfc */;
                6016: data_o = 32'h00000000 /* 0x5e00 */;
                6017: data_o = 32'h00000000 /* 0x5e04 */;
                6018: data_o = 32'h00000000 /* 0x5e08 */;
                6019: data_o = 32'h00000000 /* 0x5e0c */;
                6020: data_o = 32'h00000000 /* 0x5e10 */;
                6021: data_o = 32'h00000000 /* 0x5e14 */;
                6022: data_o = 32'h00000000 /* 0x5e18 */;
                6023: data_o = 32'h00000000 /* 0x5e1c */;
                6024: data_o = 32'h00000000 /* 0x5e20 */;
                6025: data_o = 32'h00000000 /* 0x5e24 */;
                6026: data_o = 32'h00000000 /* 0x5e28 */;
                6027: data_o = 32'h00000000 /* 0x5e2c */;
                6028: data_o = 32'h00000000 /* 0x5e30 */;
                6029: data_o = 32'h00000000 /* 0x5e34 */;
                6030: data_o = 32'h00000000 /* 0x5e38 */;
                6031: data_o = 32'h00000000 /* 0x5e3c */;
                6032: data_o = 32'h00000000 /* 0x5e40 */;
                6033: data_o = 32'h00000000 /* 0x5e44 */;
                6034: data_o = 32'h00000000 /* 0x5e48 */;
                6035: data_o = 32'h00000000 /* 0x5e4c */;
                6036: data_o = 32'h00000000 /* 0x5e50 */;
                6037: data_o = 32'h00000000 /* 0x5e54 */;
                6038: data_o = 32'h00000000 /* 0x5e58 */;
                6039: data_o = 32'h00000000 /* 0x5e5c */;
                6040: data_o = 32'h00000000 /* 0x5e60 */;
                6041: data_o = 32'h00000000 /* 0x5e64 */;
                6042: data_o = 32'h00000000 /* 0x5e68 */;
                6043: data_o = 32'h00000000 /* 0x5e6c */;
                6044: data_o = 32'h00000000 /* 0x5e70 */;
                6045: data_o = 32'h00000000 /* 0x5e74 */;
                6046: data_o = 32'h00000000 /* 0x5e78 */;
                6047: data_o = 32'h00000000 /* 0x5e7c */;
                6048: data_o = 32'h00000000 /* 0x5e80 */;
                6049: data_o = 32'h00000000 /* 0x5e84 */;
                6050: data_o = 32'h00000000 /* 0x5e88 */;
                6051: data_o = 32'h00000000 /* 0x5e8c */;
                6052: data_o = 32'h00000000 /* 0x5e90 */;
                6053: data_o = 32'h00000000 /* 0x5e94 */;
                6054: data_o = 32'h00000000 /* 0x5e98 */;
                6055: data_o = 32'h00000000 /* 0x5e9c */;
                6056: data_o = 32'h00000000 /* 0x5ea0 */;
                6057: data_o = 32'h00000000 /* 0x5ea4 */;
                6058: data_o = 32'h00000000 /* 0x5ea8 */;
                6059: data_o = 32'h00000000 /* 0x5eac */;
                6060: data_o = 32'h00000000 /* 0x5eb0 */;
                6061: data_o = 32'h00000000 /* 0x5eb4 */;
                6062: data_o = 32'h00000000 /* 0x5eb8 */;
                6063: data_o = 32'h00000000 /* 0x5ebc */;
                6064: data_o = 32'h00000000 /* 0x5ec0 */;
                6065: data_o = 32'h00000000 /* 0x5ec4 */;
                6066: data_o = 32'h00000000 /* 0x5ec8 */;
                6067: data_o = 32'h00000000 /* 0x5ecc */;
                6068: data_o = 32'h00000000 /* 0x5ed0 */;
                6069: data_o = 32'h00000000 /* 0x5ed4 */;
                6070: data_o = 32'h00000000 /* 0x5ed8 */;
                6071: data_o = 32'h00000000 /* 0x5edc */;
                6072: data_o = 32'h00000000 /* 0x5ee0 */;
                6073: data_o = 32'h00000000 /* 0x5ee4 */;
                6074: data_o = 32'h00000000 /* 0x5ee8 */;
                6075: data_o = 32'h00000000 /* 0x5eec */;
                6076: data_o = 32'h00000000 /* 0x5ef0 */;
                6077: data_o = 32'h00000000 /* 0x5ef4 */;
                6078: data_o = 32'h00000000 /* 0x5ef8 */;
                6079: data_o = 32'h00000000 /* 0x5efc */;
                6080: data_o = 32'h00000000 /* 0x5f00 */;
                6081: data_o = 32'h00000000 /* 0x5f04 */;
                6082: data_o = 32'h00000000 /* 0x5f08 */;
                6083: data_o = 32'h00000000 /* 0x5f0c */;
                6084: data_o = 32'h00000000 /* 0x5f10 */;
                6085: data_o = 32'h00000000 /* 0x5f14 */;
                6086: data_o = 32'h00000000 /* 0x5f18 */;
                6087: data_o = 32'h00000000 /* 0x5f1c */;
                6088: data_o = 32'h00000000 /* 0x5f20 */;
                6089: data_o = 32'h00000000 /* 0x5f24 */;
                6090: data_o = 32'h00000000 /* 0x5f28 */;
                6091: data_o = 32'h00000000 /* 0x5f2c */;
                6092: data_o = 32'h00000000 /* 0x5f30 */;
                6093: data_o = 32'h00000000 /* 0x5f34 */;
                6094: data_o = 32'h00000000 /* 0x5f38 */;
                6095: data_o = 32'h00000000 /* 0x5f3c */;
                6096: data_o = 32'h00000000 /* 0x5f40 */;
                6097: data_o = 32'h00000000 /* 0x5f44 */;
                6098: data_o = 32'h00000000 /* 0x5f48 */;
                6099: data_o = 32'h00000000 /* 0x5f4c */;
                6100: data_o = 32'h00000000 /* 0x5f50 */;
                6101: data_o = 32'h00000000 /* 0x5f54 */;
                6102: data_o = 32'h00000000 /* 0x5f58 */;
                6103: data_o = 32'h00000000 /* 0x5f5c */;
                6104: data_o = 32'h00000000 /* 0x5f60 */;
                6105: data_o = 32'h00000000 /* 0x5f64 */;
                6106: data_o = 32'h00000000 /* 0x5f68 */;
                6107: data_o = 32'h00000000 /* 0x5f6c */;
                6108: data_o = 32'h00000000 /* 0x5f70 */;
                6109: data_o = 32'h00000000 /* 0x5f74 */;
                6110: data_o = 32'h00000000 /* 0x5f78 */;
                6111: data_o = 32'h00000000 /* 0x5f7c */;
                6112: data_o = 32'h00000000 /* 0x5f80 */;
                6113: data_o = 32'h00000000 /* 0x5f84 */;
                6114: data_o = 32'h00000000 /* 0x5f88 */;
                6115: data_o = 32'h00000000 /* 0x5f8c */;
                6116: data_o = 32'h00000000 /* 0x5f90 */;
                6117: data_o = 32'h00000000 /* 0x5f94 */;
                6118: data_o = 32'h00000000 /* 0x5f98 */;
                6119: data_o = 32'h00000000 /* 0x5f9c */;
                6120: data_o = 32'h00000000 /* 0x5fa0 */;
                6121: data_o = 32'h00000000 /* 0x5fa4 */;
                6122: data_o = 32'h00000000 /* 0x5fa8 */;
                6123: data_o = 32'h00000000 /* 0x5fac */;
                6124: data_o = 32'h00000000 /* 0x5fb0 */;
                6125: data_o = 32'h00000000 /* 0x5fb4 */;
                6126: data_o = 32'h00000000 /* 0x5fb8 */;
                6127: data_o = 32'h00000000 /* 0x5fbc */;
                6128: data_o = 32'h00000000 /* 0x5fc0 */;
                6129: data_o = 32'h00000000 /* 0x5fc4 */;
                6130: data_o = 32'h00000000 /* 0x5fc8 */;
                6131: data_o = 32'h00000000 /* 0x5fcc */;
                6132: data_o = 32'h00000000 /* 0x5fd0 */;
                6133: data_o = 32'h00000000 /* 0x5fd4 */;
                6134: data_o = 32'h00000000 /* 0x5fd8 */;
                6135: data_o = 32'h00000000 /* 0x5fdc */;
                6136: data_o = 32'h00000000 /* 0x5fe0 */;
                6137: data_o = 32'h00000000 /* 0x5fe4 */;
                6138: data_o = 32'h00000000 /* 0x5fe8 */;
                6139: data_o = 32'h00000000 /* 0x5fec */;
                6140: data_o = 32'h00000000 /* 0x5ff0 */;
                6141: data_o = 32'h00000000 /* 0x5ff4 */;
                6142: data_o = 32'h00000000 /* 0x5ff8 */;
                6143: data_o = 32'h00000000 /* 0x5ffc */;
                6144: data_o = 32'h00000000 /* 0x6000 */;
                6145: data_o = 32'h00000000 /* 0x6004 */;
                6146: data_o = 32'h00000000 /* 0x6008 */;
                6147: data_o = 32'h00000000 /* 0x600c */;
                6148: data_o = 32'h00000000 /* 0x6010 */;
                6149: data_o = 32'h00000000 /* 0x6014 */;
                6150: data_o = 32'h00000000 /* 0x6018 */;
                6151: data_o = 32'h00000000 /* 0x601c */;
                6152: data_o = 32'h00000000 /* 0x6020 */;
                6153: data_o = 32'h00000000 /* 0x6024 */;
                6154: data_o = 32'h00000000 /* 0x6028 */;
                6155: data_o = 32'h00000000 /* 0x602c */;
                6156: data_o = 32'h00000000 /* 0x6030 */;
                6157: data_o = 32'h00000000 /* 0x6034 */;
                6158: data_o = 32'h00000000 /* 0x6038 */;
                6159: data_o = 32'h00000000 /* 0x603c */;
                6160: data_o = 32'h00000000 /* 0x6040 */;
                6161: data_o = 32'h00000000 /* 0x6044 */;
                6162: data_o = 32'h00000000 /* 0x6048 */;
                6163: data_o = 32'h00000000 /* 0x604c */;
                6164: data_o = 32'h00000000 /* 0x6050 */;
                6165: data_o = 32'h00000000 /* 0x6054 */;
                6166: data_o = 32'h00000000 /* 0x6058 */;
                6167: data_o = 32'h00000000 /* 0x605c */;
                6168: data_o = 32'h00000000 /* 0x6060 */;
                6169: data_o = 32'h00000000 /* 0x6064 */;
                6170: data_o = 32'h00000000 /* 0x6068 */;
                6171: data_o = 32'h00000000 /* 0x606c */;
                6172: data_o = 32'h00000000 /* 0x6070 */;
                6173: data_o = 32'h00000000 /* 0x6074 */;
                6174: data_o = 32'h00000000 /* 0x6078 */;
                6175: data_o = 32'h00000000 /* 0x607c */;
                6176: data_o = 32'h00000000 /* 0x6080 */;
                6177: data_o = 32'h00000000 /* 0x6084 */;
                6178: data_o = 32'h00000000 /* 0x6088 */;
                6179: data_o = 32'h00000000 /* 0x608c */;
                6180: data_o = 32'h00000000 /* 0x6090 */;
                6181: data_o = 32'h00000000 /* 0x6094 */;
                6182: data_o = 32'h00000000 /* 0x6098 */;
                6183: data_o = 32'h00000000 /* 0x609c */;
                6184: data_o = 32'h00000000 /* 0x60a0 */;
                6185: data_o = 32'h00000000 /* 0x60a4 */;
                6186: data_o = 32'h00000000 /* 0x60a8 */;
                6187: data_o = 32'h00000000 /* 0x60ac */;
                6188: data_o = 32'h00000000 /* 0x60b0 */;
                6189: data_o = 32'h00000000 /* 0x60b4 */;
                6190: data_o = 32'h00000000 /* 0x60b8 */;
                6191: data_o = 32'h00000000 /* 0x60bc */;
                6192: data_o = 32'h00000000 /* 0x60c0 */;
                6193: data_o = 32'h00000000 /* 0x60c4 */;
                6194: data_o = 32'h00000000 /* 0x60c8 */;
                6195: data_o = 32'h00000000 /* 0x60cc */;
                6196: data_o = 32'h00000000 /* 0x60d0 */;
                6197: data_o = 32'h00000000 /* 0x60d4 */;
                6198: data_o = 32'h00000000 /* 0x60d8 */;
                6199: data_o = 32'h00000000 /* 0x60dc */;
                6200: data_o = 32'h00000000 /* 0x60e0 */;
                6201: data_o = 32'h00000000 /* 0x60e4 */;
                6202: data_o = 32'h00000000 /* 0x60e8 */;
                6203: data_o = 32'h00000000 /* 0x60ec */;
                6204: data_o = 32'h00000000 /* 0x60f0 */;
                6205: data_o = 32'h00000000 /* 0x60f4 */;
                6206: data_o = 32'h00000000 /* 0x60f8 */;
                6207: data_o = 32'h00000000 /* 0x60fc */;
                6208: data_o = 32'h00000000 /* 0x6100 */;
                6209: data_o = 32'h00000000 /* 0x6104 */;
                6210: data_o = 32'h00000000 /* 0x6108 */;
                6211: data_o = 32'h00000000 /* 0x610c */;
                6212: data_o = 32'h00000000 /* 0x6110 */;
                6213: data_o = 32'h00000000 /* 0x6114 */;
                6214: data_o = 32'h00000000 /* 0x6118 */;
                6215: data_o = 32'h00000000 /* 0x611c */;
                6216: data_o = 32'h00000000 /* 0x6120 */;
                6217: data_o = 32'h00000000 /* 0x6124 */;
                6218: data_o = 32'h00000000 /* 0x6128 */;
                6219: data_o = 32'h00000000 /* 0x612c */;
                6220: data_o = 32'h00000000 /* 0x6130 */;
                6221: data_o = 32'h00000000 /* 0x6134 */;
                6222: data_o = 32'h00000000 /* 0x6138 */;
                6223: data_o = 32'h00000000 /* 0x613c */;
                6224: data_o = 32'h00000000 /* 0x6140 */;
                6225: data_o = 32'h00000000 /* 0x6144 */;
                6226: data_o = 32'h00000000 /* 0x6148 */;
                6227: data_o = 32'h00000000 /* 0x614c */;
                6228: data_o = 32'h00000000 /* 0x6150 */;
                6229: data_o = 32'h00000000 /* 0x6154 */;
                6230: data_o = 32'h00000000 /* 0x6158 */;
                6231: data_o = 32'h00000000 /* 0x615c */;
                6232: data_o = 32'h00000000 /* 0x6160 */;
                6233: data_o = 32'h00000000 /* 0x6164 */;
                6234: data_o = 32'h00000000 /* 0x6168 */;
                6235: data_o = 32'h00000000 /* 0x616c */;
                6236: data_o = 32'h00000000 /* 0x6170 */;
                6237: data_o = 32'h00000000 /* 0x6174 */;
                6238: data_o = 32'h00000000 /* 0x6178 */;
                6239: data_o = 32'h00000000 /* 0x617c */;
                6240: data_o = 32'h00000000 /* 0x6180 */;
                6241: data_o = 32'h00000000 /* 0x6184 */;
                6242: data_o = 32'h00000000 /* 0x6188 */;
                6243: data_o = 32'h00000000 /* 0x618c */;
                6244: data_o = 32'h00000000 /* 0x6190 */;
                6245: data_o = 32'h00000000 /* 0x6194 */;
                6246: data_o = 32'h00000000 /* 0x6198 */;
                6247: data_o = 32'h00000000 /* 0x619c */;
                6248: data_o = 32'h00000000 /* 0x61a0 */;
                6249: data_o = 32'h00000000 /* 0x61a4 */;
                6250: data_o = 32'h00000000 /* 0x61a8 */;
                6251: data_o = 32'h00000000 /* 0x61ac */;
                6252: data_o = 32'h00000000 /* 0x61b0 */;
                6253: data_o = 32'h00000000 /* 0x61b4 */;
                6254: data_o = 32'h00000000 /* 0x61b8 */;
                6255: data_o = 32'h00000000 /* 0x61bc */;
                6256: data_o = 32'h00000000 /* 0x61c0 */;
                6257: data_o = 32'h00000000 /* 0x61c4 */;
                6258: data_o = 32'h00000000 /* 0x61c8 */;
                6259: data_o = 32'h00000000 /* 0x61cc */;
                6260: data_o = 32'h00000000 /* 0x61d0 */;
                6261: data_o = 32'h00000000 /* 0x61d4 */;
                6262: data_o = 32'h00000000 /* 0x61d8 */;
                6263: data_o = 32'h00000000 /* 0x61dc */;
                6264: data_o = 32'h00000000 /* 0x61e0 */;
                6265: data_o = 32'h00000000 /* 0x61e4 */;
                6266: data_o = 32'h00000000 /* 0x61e8 */;
                6267: data_o = 32'h00000000 /* 0x61ec */;
                6268: data_o = 32'h00000000 /* 0x61f0 */;
                6269: data_o = 32'h00000000 /* 0x61f4 */;
                6270: data_o = 32'h00000000 /* 0x61f8 */;
                6271: data_o = 32'h00000000 /* 0x61fc */;
                6272: data_o = 32'h00000000 /* 0x6200 */;
                6273: data_o = 32'h00000000 /* 0x6204 */;
                6274: data_o = 32'h00000000 /* 0x6208 */;
                6275: data_o = 32'h00000000 /* 0x620c */;
                6276: data_o = 32'h00000000 /* 0x6210 */;
                6277: data_o = 32'h00000000 /* 0x6214 */;
                6278: data_o = 32'h00000000 /* 0x6218 */;
                6279: data_o = 32'h00000000 /* 0x621c */;
                6280: data_o = 32'h00000000 /* 0x6220 */;
                6281: data_o = 32'h00000000 /* 0x6224 */;
                6282: data_o = 32'h00000000 /* 0x6228 */;
                6283: data_o = 32'h00000000 /* 0x622c */;
                6284: data_o = 32'h00000000 /* 0x6230 */;
                6285: data_o = 32'h00000000 /* 0x6234 */;
                6286: data_o = 32'h00000000 /* 0x6238 */;
                6287: data_o = 32'h00000000 /* 0x623c */;
                6288: data_o = 32'h00000000 /* 0x6240 */;
                6289: data_o = 32'h00000000 /* 0x6244 */;
                6290: data_o = 32'h00000000 /* 0x6248 */;
                6291: data_o = 32'h00000000 /* 0x624c */;
                6292: data_o = 32'h00000000 /* 0x6250 */;
                6293: data_o = 32'h00000000 /* 0x6254 */;
                6294: data_o = 32'h00000000 /* 0x6258 */;
                6295: data_o = 32'h00000000 /* 0x625c */;
                6296: data_o = 32'h00000000 /* 0x6260 */;
                6297: data_o = 32'h00000000 /* 0x6264 */;
                6298: data_o = 32'h00000000 /* 0x6268 */;
                6299: data_o = 32'h00000000 /* 0x626c */;
                6300: data_o = 32'h00000000 /* 0x6270 */;
                6301: data_o = 32'h00000000 /* 0x6274 */;
                6302: data_o = 32'h00000000 /* 0x6278 */;
                6303: data_o = 32'h00000000 /* 0x627c */;
                6304: data_o = 32'h00000000 /* 0x6280 */;
                6305: data_o = 32'h00000000 /* 0x6284 */;
                6306: data_o = 32'h00000000 /* 0x6288 */;
                6307: data_o = 32'h00000000 /* 0x628c */;
                6308: data_o = 32'h00000000 /* 0x6290 */;
                6309: data_o = 32'h00000000 /* 0x6294 */;
                6310: data_o = 32'h00000000 /* 0x6298 */;
                6311: data_o = 32'h00000000 /* 0x629c */;
                6312: data_o = 32'h00000000 /* 0x62a0 */;
                6313: data_o = 32'h00000000 /* 0x62a4 */;
                6314: data_o = 32'h00000000 /* 0x62a8 */;
                6315: data_o = 32'h00000000 /* 0x62ac */;
                6316: data_o = 32'h00000000 /* 0x62b0 */;
                6317: data_o = 32'h00000000 /* 0x62b4 */;
                6318: data_o = 32'h00000000 /* 0x62b8 */;
                6319: data_o = 32'h00000000 /* 0x62bc */;
                6320: data_o = 32'h00000000 /* 0x62c0 */;
                6321: data_o = 32'h00000000 /* 0x62c4 */;
                6322: data_o = 32'h00000000 /* 0x62c8 */;
                6323: data_o = 32'h00000000 /* 0x62cc */;
                6324: data_o = 32'h00000000 /* 0x62d0 */;
                6325: data_o = 32'h00000000 /* 0x62d4 */;
                6326: data_o = 32'h00000000 /* 0x62d8 */;
                6327: data_o = 32'h00000000 /* 0x62dc */;
                6328: data_o = 32'h00000000 /* 0x62e0 */;
                6329: data_o = 32'h00000000 /* 0x62e4 */;
                6330: data_o = 32'h00000000 /* 0x62e8 */;
                6331: data_o = 32'h00000000 /* 0x62ec */;
                6332: data_o = 32'h00000000 /* 0x62f0 */;
                6333: data_o = 32'h00000000 /* 0x62f4 */;
                6334: data_o = 32'h00000000 /* 0x62f8 */;
                6335: data_o = 32'h00000000 /* 0x62fc */;
                6336: data_o = 32'h00000000 /* 0x6300 */;
                6337: data_o = 32'h00000000 /* 0x6304 */;
                6338: data_o = 32'h00000000 /* 0x6308 */;
                6339: data_o = 32'h00000000 /* 0x630c */;
                6340: data_o = 32'h00000000 /* 0x6310 */;
                6341: data_o = 32'h00000000 /* 0x6314 */;
                6342: data_o = 32'h00000000 /* 0x6318 */;
                6343: data_o = 32'h00000000 /* 0x631c */;
                6344: data_o = 32'h00000000 /* 0x6320 */;
                6345: data_o = 32'h00000000 /* 0x6324 */;
                6346: data_o = 32'h00000000 /* 0x6328 */;
                6347: data_o = 32'h00000000 /* 0x632c */;
                6348: data_o = 32'h00000000 /* 0x6330 */;
                6349: data_o = 32'h00000000 /* 0x6334 */;
                6350: data_o = 32'h00000000 /* 0x6338 */;
                6351: data_o = 32'h00000000 /* 0x633c */;
                6352: data_o = 32'h00000000 /* 0x6340 */;
                6353: data_o = 32'h00000000 /* 0x6344 */;
                6354: data_o = 32'h00000000 /* 0x6348 */;
                6355: data_o = 32'h00000000 /* 0x634c */;
                6356: data_o = 32'h00000000 /* 0x6350 */;
                6357: data_o = 32'h00000000 /* 0x6354 */;
                6358: data_o = 32'h00000000 /* 0x6358 */;
                6359: data_o = 32'h00000000 /* 0x635c */;
                6360: data_o = 32'h00000000 /* 0x6360 */;
                6361: data_o = 32'h00000000 /* 0x6364 */;
                6362: data_o = 32'h00000000 /* 0x6368 */;
                6363: data_o = 32'h00000000 /* 0x636c */;
                6364: data_o = 32'h00000000 /* 0x6370 */;
                6365: data_o = 32'h00000000 /* 0x6374 */;
                6366: data_o = 32'h00000000 /* 0x6378 */;
                6367: data_o = 32'h00000000 /* 0x637c */;
                6368: data_o = 32'h00000000 /* 0x6380 */;
                6369: data_o = 32'h00000000 /* 0x6384 */;
                6370: data_o = 32'h00000000 /* 0x6388 */;
                6371: data_o = 32'h00000000 /* 0x638c */;
                6372: data_o = 32'h00000000 /* 0x6390 */;
                6373: data_o = 32'h00000000 /* 0x6394 */;
                6374: data_o = 32'h00000000 /* 0x6398 */;
                6375: data_o = 32'h00000000 /* 0x639c */;
                6376: data_o = 32'h00000000 /* 0x63a0 */;
                6377: data_o = 32'h00000000 /* 0x63a4 */;
                6378: data_o = 32'h00000000 /* 0x63a8 */;
                6379: data_o = 32'h00000000 /* 0x63ac */;
                6380: data_o = 32'h00000000 /* 0x63b0 */;
                6381: data_o = 32'h00000000 /* 0x63b4 */;
                6382: data_o = 32'h00000000 /* 0x63b8 */;
                6383: data_o = 32'h00000000 /* 0x63bc */;
                6384: data_o = 32'h00000000 /* 0x63c0 */;
                6385: data_o = 32'h00000000 /* 0x63c4 */;
                6386: data_o = 32'h00000000 /* 0x63c8 */;
                6387: data_o = 32'h00000000 /* 0x63cc */;
                6388: data_o = 32'h00000000 /* 0x63d0 */;
                6389: data_o = 32'h00000000 /* 0x63d4 */;
                6390: data_o = 32'h00000000 /* 0x63d8 */;
                6391: data_o = 32'h00000000 /* 0x63dc */;
                6392: data_o = 32'h00000000 /* 0x63e0 */;
                6393: data_o = 32'h00000000 /* 0x63e4 */;
                6394: data_o = 32'h00000000 /* 0x63e8 */;
                6395: data_o = 32'h00000000 /* 0x63ec */;
                6396: data_o = 32'h00000000 /* 0x63f0 */;
                6397: data_o = 32'h00000000 /* 0x63f4 */;
                6398: data_o = 32'h00000000 /* 0x63f8 */;
                6399: data_o = 32'h00000000 /* 0x63fc */;
                6400: data_o = 32'h00000000 /* 0x6400 */;
                6401: data_o = 32'h00000000 /* 0x6404 */;
                6402: data_o = 32'h00000000 /* 0x6408 */;
                6403: data_o = 32'h00000000 /* 0x640c */;
                6404: data_o = 32'h00000000 /* 0x6410 */;
                6405: data_o = 32'h00000000 /* 0x6414 */;
                6406: data_o = 32'h00000000 /* 0x6418 */;
                6407: data_o = 32'h00000000 /* 0x641c */;
                6408: data_o = 32'h00000000 /* 0x6420 */;
                6409: data_o = 32'h00000000 /* 0x6424 */;
                6410: data_o = 32'h00000000 /* 0x6428 */;
                6411: data_o = 32'h00000000 /* 0x642c */;
                6412: data_o = 32'h00000000 /* 0x6430 */;
                6413: data_o = 32'h00000000 /* 0x6434 */;
                6414: data_o = 32'h00000000 /* 0x6438 */;
                6415: data_o = 32'h00000000 /* 0x643c */;
                6416: data_o = 32'h00000000 /* 0x6440 */;
                6417: data_o = 32'h00000000 /* 0x6444 */;
                6418: data_o = 32'h00000000 /* 0x6448 */;
                6419: data_o = 32'h00000000 /* 0x644c */;
                6420: data_o = 32'h00000000 /* 0x6450 */;
                6421: data_o = 32'h00000000 /* 0x6454 */;
                6422: data_o = 32'h00000000 /* 0x6458 */;
                6423: data_o = 32'h00000000 /* 0x645c */;
                6424: data_o = 32'h00000000 /* 0x6460 */;
                6425: data_o = 32'h00000000 /* 0x6464 */;
                6426: data_o = 32'h00000000 /* 0x6468 */;
                6427: data_o = 32'h00000000 /* 0x646c */;
                6428: data_o = 32'h00000000 /* 0x6470 */;
                6429: data_o = 32'h00000000 /* 0x6474 */;
                6430: data_o = 32'h00000000 /* 0x6478 */;
                6431: data_o = 32'h00000000 /* 0x647c */;
                6432: data_o = 32'h00000000 /* 0x6480 */;
                6433: data_o = 32'h00000000 /* 0x6484 */;
                6434: data_o = 32'h00000000 /* 0x6488 */;
                6435: data_o = 32'h00000000 /* 0x648c */;
                6436: data_o = 32'h00000000 /* 0x6490 */;
                6437: data_o = 32'h00000000 /* 0x6494 */;
                6438: data_o = 32'h00000000 /* 0x6498 */;
                6439: data_o = 32'h00000000 /* 0x649c */;
                6440: data_o = 32'h00000000 /* 0x64a0 */;
                6441: data_o = 32'h00000000 /* 0x64a4 */;
                6442: data_o = 32'h00000000 /* 0x64a8 */;
                6443: data_o = 32'h00000000 /* 0x64ac */;
                6444: data_o = 32'h00000000 /* 0x64b0 */;
                6445: data_o = 32'h00000000 /* 0x64b4 */;
                6446: data_o = 32'h00000000 /* 0x64b8 */;
                6447: data_o = 32'h00000000 /* 0x64bc */;
                6448: data_o = 32'h00000000 /* 0x64c0 */;
                6449: data_o = 32'h00000000 /* 0x64c4 */;
                6450: data_o = 32'h00000000 /* 0x64c8 */;
                6451: data_o = 32'h00000000 /* 0x64cc */;
                6452: data_o = 32'h00000000 /* 0x64d0 */;
                6453: data_o = 32'h00000000 /* 0x64d4 */;
                6454: data_o = 32'h00000000 /* 0x64d8 */;
                6455: data_o = 32'h00000000 /* 0x64dc */;
                6456: data_o = 32'h00000000 /* 0x64e0 */;
                6457: data_o = 32'h00000000 /* 0x64e4 */;
                6458: data_o = 32'h00000000 /* 0x64e8 */;
                6459: data_o = 32'h00000000 /* 0x64ec */;
                6460: data_o = 32'h00000000 /* 0x64f0 */;
                6461: data_o = 32'h00000000 /* 0x64f4 */;
                6462: data_o = 32'h00000000 /* 0x64f8 */;
                6463: data_o = 32'h00000000 /* 0x64fc */;
                6464: data_o = 32'h00000000 /* 0x6500 */;
                6465: data_o = 32'h00000000 /* 0x6504 */;
                6466: data_o = 32'h00000000 /* 0x6508 */;
                6467: data_o = 32'h00000000 /* 0x650c */;
                6468: data_o = 32'h00000000 /* 0x6510 */;
                6469: data_o = 32'h00000000 /* 0x6514 */;
                6470: data_o = 32'h00000000 /* 0x6518 */;
                6471: data_o = 32'h00000000 /* 0x651c */;
                6472: data_o = 32'h00000000 /* 0x6520 */;
                6473: data_o = 32'h00000000 /* 0x6524 */;
                6474: data_o = 32'h00000000 /* 0x6528 */;
                6475: data_o = 32'h00000000 /* 0x652c */;
                6476: data_o = 32'h00000000 /* 0x6530 */;
                6477: data_o = 32'h00000000 /* 0x6534 */;
                6478: data_o = 32'h00000000 /* 0x6538 */;
                6479: data_o = 32'h00000000 /* 0x653c */;
                6480: data_o = 32'h00000000 /* 0x6540 */;
                6481: data_o = 32'h00000000 /* 0x6544 */;
                6482: data_o = 32'h00000000 /* 0x6548 */;
                6483: data_o = 32'h00000000 /* 0x654c */;
                6484: data_o = 32'h00000000 /* 0x6550 */;
                6485: data_o = 32'h00000000 /* 0x6554 */;
                6486: data_o = 32'h00000000 /* 0x6558 */;
                6487: data_o = 32'h00000000 /* 0x655c */;
                6488: data_o = 32'h00000000 /* 0x6560 */;
                6489: data_o = 32'h00000000 /* 0x6564 */;
                6490: data_o = 32'h00000000 /* 0x6568 */;
                6491: data_o = 32'h00000000 /* 0x656c */;
                6492: data_o = 32'h00000000 /* 0x6570 */;
                6493: data_o = 32'h00000000 /* 0x6574 */;
                6494: data_o = 32'h00000000 /* 0x6578 */;
                6495: data_o = 32'h00000000 /* 0x657c */;
                6496: data_o = 32'h00000000 /* 0x6580 */;
                6497: data_o = 32'h00000000 /* 0x6584 */;
                6498: data_o = 32'h00000000 /* 0x6588 */;
                6499: data_o = 32'h00000000 /* 0x658c */;
                6500: data_o = 32'h00000000 /* 0x6590 */;
                6501: data_o = 32'h00000000 /* 0x6594 */;
                6502: data_o = 32'h00000000 /* 0x6598 */;
                6503: data_o = 32'h00000000 /* 0x659c */;
                6504: data_o = 32'h00000000 /* 0x65a0 */;
                6505: data_o = 32'h00000000 /* 0x65a4 */;
                6506: data_o = 32'h00000000 /* 0x65a8 */;
                6507: data_o = 32'h00000000 /* 0x65ac */;
                6508: data_o = 32'h00000000 /* 0x65b0 */;
                6509: data_o = 32'h00000000 /* 0x65b4 */;
                6510: data_o = 32'h00000000 /* 0x65b8 */;
                6511: data_o = 32'h00000000 /* 0x65bc */;
                6512: data_o = 32'h00000000 /* 0x65c0 */;
                6513: data_o = 32'h00000000 /* 0x65c4 */;
                6514: data_o = 32'h00000000 /* 0x65c8 */;
                6515: data_o = 32'h00000000 /* 0x65cc */;
                6516: data_o = 32'h00000000 /* 0x65d0 */;
                6517: data_o = 32'h00000000 /* 0x65d4 */;
                6518: data_o = 32'h00000000 /* 0x65d8 */;
                6519: data_o = 32'h00000000 /* 0x65dc */;
                6520: data_o = 32'h00000000 /* 0x65e0 */;
                6521: data_o = 32'h00000000 /* 0x65e4 */;
                6522: data_o = 32'h00000000 /* 0x65e8 */;
                6523: data_o = 32'h00000000 /* 0x65ec */;
                6524: data_o = 32'h00000000 /* 0x65f0 */;
                6525: data_o = 32'h00000000 /* 0x65f4 */;
                6526: data_o = 32'h00000000 /* 0x65f8 */;
                6527: data_o = 32'h00000000 /* 0x65fc */;
                6528: data_o = 32'h00000000 /* 0x6600 */;
                6529: data_o = 32'h00000000 /* 0x6604 */;
                6530: data_o = 32'h00000000 /* 0x6608 */;
                6531: data_o = 32'h00000000 /* 0x660c */;
                6532: data_o = 32'h00000000 /* 0x6610 */;
                6533: data_o = 32'h00000000 /* 0x6614 */;
                6534: data_o = 32'h00000000 /* 0x6618 */;
                6535: data_o = 32'h00000000 /* 0x661c */;
                6536: data_o = 32'h00000000 /* 0x6620 */;
                6537: data_o = 32'h00000000 /* 0x6624 */;
                6538: data_o = 32'h00000000 /* 0x6628 */;
                6539: data_o = 32'h00000000 /* 0x662c */;
                6540: data_o = 32'h00000000 /* 0x6630 */;
                6541: data_o = 32'h00000000 /* 0x6634 */;
                6542: data_o = 32'h00000000 /* 0x6638 */;
                6543: data_o = 32'h00000000 /* 0x663c */;
                6544: data_o = 32'h00000000 /* 0x6640 */;
                6545: data_o = 32'h00000000 /* 0x6644 */;
                6546: data_o = 32'h00000000 /* 0x6648 */;
                6547: data_o = 32'h00000000 /* 0x664c */;
                6548: data_o = 32'h00000000 /* 0x6650 */;
                6549: data_o = 32'h00000000 /* 0x6654 */;
                6550: data_o = 32'h00000000 /* 0x6658 */;
                6551: data_o = 32'h00000000 /* 0x665c */;
                6552: data_o = 32'h00000000 /* 0x6660 */;
                6553: data_o = 32'h00000000 /* 0x6664 */;
                6554: data_o = 32'h00000000 /* 0x6668 */;
                6555: data_o = 32'h00000000 /* 0x666c */;
                6556: data_o = 32'h00000000 /* 0x6670 */;
                6557: data_o = 32'h00000000 /* 0x6674 */;
                6558: data_o = 32'h00000000 /* 0x6678 */;
                6559: data_o = 32'h00000000 /* 0x667c */;
                6560: data_o = 32'h00000000 /* 0x6680 */;
                6561: data_o = 32'h00000000 /* 0x6684 */;
                6562: data_o = 32'h00000000 /* 0x6688 */;
                6563: data_o = 32'h00000000 /* 0x668c */;
                6564: data_o = 32'h00000000 /* 0x6690 */;
                6565: data_o = 32'h00000000 /* 0x6694 */;
                6566: data_o = 32'h00000000 /* 0x6698 */;
                6567: data_o = 32'h00000000 /* 0x669c */;
                6568: data_o = 32'h00000000 /* 0x66a0 */;
                6569: data_o = 32'h00000000 /* 0x66a4 */;
                6570: data_o = 32'h00000000 /* 0x66a8 */;
                6571: data_o = 32'h00000000 /* 0x66ac */;
                6572: data_o = 32'h00000000 /* 0x66b0 */;
                6573: data_o = 32'h00000000 /* 0x66b4 */;
                6574: data_o = 32'h00000000 /* 0x66b8 */;
                6575: data_o = 32'h00000000 /* 0x66bc */;
                6576: data_o = 32'h00000000 /* 0x66c0 */;
                6577: data_o = 32'h00000000 /* 0x66c4 */;
                6578: data_o = 32'h00000000 /* 0x66c8 */;
                6579: data_o = 32'h00000000 /* 0x66cc */;
                6580: data_o = 32'h00000000 /* 0x66d0 */;
                6581: data_o = 32'h00000000 /* 0x66d4 */;
                6582: data_o = 32'h00000000 /* 0x66d8 */;
                6583: data_o = 32'h00000000 /* 0x66dc */;
                6584: data_o = 32'h00000000 /* 0x66e0 */;
                6585: data_o = 32'h00000000 /* 0x66e4 */;
                6586: data_o = 32'h00000000 /* 0x66e8 */;
                6587: data_o = 32'h00000000 /* 0x66ec */;
                6588: data_o = 32'h00000000 /* 0x66f0 */;
                6589: data_o = 32'h00000000 /* 0x66f4 */;
                6590: data_o = 32'h00000000 /* 0x66f8 */;
                6591: data_o = 32'h00000000 /* 0x66fc */;
                6592: data_o = 32'h00000000 /* 0x6700 */;
                6593: data_o = 32'h00000000 /* 0x6704 */;
                6594: data_o = 32'h00000000 /* 0x6708 */;
                6595: data_o = 32'h00000000 /* 0x670c */;
                6596: data_o = 32'h00000000 /* 0x6710 */;
                6597: data_o = 32'h00000000 /* 0x6714 */;
                6598: data_o = 32'h00000000 /* 0x6718 */;
                6599: data_o = 32'h00000000 /* 0x671c */;
                6600: data_o = 32'h00000000 /* 0x6720 */;
                6601: data_o = 32'h00000000 /* 0x6724 */;
                6602: data_o = 32'h00000000 /* 0x6728 */;
                6603: data_o = 32'h00000000 /* 0x672c */;
                6604: data_o = 32'h00000000 /* 0x6730 */;
                6605: data_o = 32'h00000000 /* 0x6734 */;
                6606: data_o = 32'h00000000 /* 0x6738 */;
                6607: data_o = 32'h00000000 /* 0x673c */;
                6608: data_o = 32'h00000000 /* 0x6740 */;
                6609: data_o = 32'h00000000 /* 0x6744 */;
                6610: data_o = 32'h00000000 /* 0x6748 */;
                6611: data_o = 32'h00000000 /* 0x674c */;
                6612: data_o = 32'h00000000 /* 0x6750 */;
                6613: data_o = 32'h00000000 /* 0x6754 */;
                6614: data_o = 32'h00000000 /* 0x6758 */;
                6615: data_o = 32'h00000000 /* 0x675c */;
                6616: data_o = 32'h00000000 /* 0x6760 */;
                6617: data_o = 32'h00000000 /* 0x6764 */;
                6618: data_o = 32'h00000000 /* 0x6768 */;
                6619: data_o = 32'h00000000 /* 0x676c */;
                6620: data_o = 32'h00000000 /* 0x6770 */;
                6621: data_o = 32'h00000000 /* 0x6774 */;
                6622: data_o = 32'h00000000 /* 0x6778 */;
                6623: data_o = 32'h00000000 /* 0x677c */;
                6624: data_o = 32'h00000000 /* 0x6780 */;
                6625: data_o = 32'h00000000 /* 0x6784 */;
                6626: data_o = 32'h00000000 /* 0x6788 */;
                6627: data_o = 32'h00000000 /* 0x678c */;
                6628: data_o = 32'h00000000 /* 0x6790 */;
                6629: data_o = 32'h00000000 /* 0x6794 */;
                6630: data_o = 32'h00000000 /* 0x6798 */;
                6631: data_o = 32'h00000000 /* 0x679c */;
                6632: data_o = 32'h00000000 /* 0x67a0 */;
                6633: data_o = 32'h00000000 /* 0x67a4 */;
                6634: data_o = 32'h00000000 /* 0x67a8 */;
                6635: data_o = 32'h00000000 /* 0x67ac */;
                6636: data_o = 32'h00000000 /* 0x67b0 */;
                6637: data_o = 32'h00000000 /* 0x67b4 */;
                6638: data_o = 32'h00000000 /* 0x67b8 */;
                6639: data_o = 32'h00000000 /* 0x67bc */;
                6640: data_o = 32'h00000000 /* 0x67c0 */;
                6641: data_o = 32'h00000000 /* 0x67c4 */;
                6642: data_o = 32'h00000000 /* 0x67c8 */;
                6643: data_o = 32'h00000000 /* 0x67cc */;
                6644: data_o = 32'h00000000 /* 0x67d0 */;
                6645: data_o = 32'h00000000 /* 0x67d4 */;
                6646: data_o = 32'h00000000 /* 0x67d8 */;
                6647: data_o = 32'h00000000 /* 0x67dc */;
                6648: data_o = 32'h00000000 /* 0x67e0 */;
                6649: data_o = 32'h00000000 /* 0x67e4 */;
                6650: data_o = 32'h00000000 /* 0x67e8 */;
                6651: data_o = 32'h00000000 /* 0x67ec */;
                6652: data_o = 32'h00000000 /* 0x67f0 */;
                6653: data_o = 32'h00000000 /* 0x67f4 */;
                6654: data_o = 32'h00000000 /* 0x67f8 */;
                6655: data_o = 32'h00000000 /* 0x67fc */;
                6656: data_o = 32'h00000000 /* 0x6800 */;
                6657: data_o = 32'h00000000 /* 0x6804 */;
                6658: data_o = 32'h00000000 /* 0x6808 */;
                6659: data_o = 32'h00000000 /* 0x680c */;
                6660: data_o = 32'h00000000 /* 0x6810 */;
                6661: data_o = 32'h00000000 /* 0x6814 */;
                6662: data_o = 32'h00000000 /* 0x6818 */;
                6663: data_o = 32'h00000000 /* 0x681c */;
                6664: data_o = 32'h00000000 /* 0x6820 */;
                6665: data_o = 32'h00000000 /* 0x6824 */;
                6666: data_o = 32'h00000000 /* 0x6828 */;
                6667: data_o = 32'h00000000 /* 0x682c */;
                6668: data_o = 32'h00000000 /* 0x6830 */;
                6669: data_o = 32'h00000000 /* 0x6834 */;
                6670: data_o = 32'h00000000 /* 0x6838 */;
                6671: data_o = 32'h00000000 /* 0x683c */;
                6672: data_o = 32'h00000000 /* 0x6840 */;
                6673: data_o = 32'h00000000 /* 0x6844 */;
                6674: data_o = 32'h00000000 /* 0x6848 */;
                6675: data_o = 32'h00000000 /* 0x684c */;
                6676: data_o = 32'h00000000 /* 0x6850 */;
                6677: data_o = 32'h00000000 /* 0x6854 */;
                6678: data_o = 32'h00000000 /* 0x6858 */;
                6679: data_o = 32'h00000000 /* 0x685c */;
                6680: data_o = 32'h00000000 /* 0x6860 */;
                6681: data_o = 32'h00000000 /* 0x6864 */;
                6682: data_o = 32'h00000000 /* 0x6868 */;
                6683: data_o = 32'h00000000 /* 0x686c */;
                6684: data_o = 32'h00000000 /* 0x6870 */;
                6685: data_o = 32'h00000000 /* 0x6874 */;
                6686: data_o = 32'h00000000 /* 0x6878 */;
                6687: data_o = 32'h00000000 /* 0x687c */;
                6688: data_o = 32'h00000000 /* 0x6880 */;
                6689: data_o = 32'h00000000 /* 0x6884 */;
                6690: data_o = 32'h00000000 /* 0x6888 */;
                6691: data_o = 32'h00000000 /* 0x688c */;
                6692: data_o = 32'h00000000 /* 0x6890 */;
                6693: data_o = 32'h00000000 /* 0x6894 */;
                6694: data_o = 32'h00000000 /* 0x6898 */;
                6695: data_o = 32'h00000000 /* 0x689c */;
                6696: data_o = 32'h00000000 /* 0x68a0 */;
                6697: data_o = 32'h00000000 /* 0x68a4 */;
                6698: data_o = 32'h00000000 /* 0x68a8 */;
                6699: data_o = 32'h00000000 /* 0x68ac */;
                6700: data_o = 32'h00000000 /* 0x68b0 */;
                6701: data_o = 32'h00000000 /* 0x68b4 */;
                6702: data_o = 32'h00000000 /* 0x68b8 */;
                6703: data_o = 32'h00000000 /* 0x68bc */;
                6704: data_o = 32'h00000000 /* 0x68c0 */;
                6705: data_o = 32'h00000000 /* 0x68c4 */;
                6706: data_o = 32'h00000000 /* 0x68c8 */;
                6707: data_o = 32'h00000000 /* 0x68cc */;
                6708: data_o = 32'h00000000 /* 0x68d0 */;
                6709: data_o = 32'h00000000 /* 0x68d4 */;
                6710: data_o = 32'h00000000 /* 0x68d8 */;
                6711: data_o = 32'h00000000 /* 0x68dc */;
                6712: data_o = 32'h00000000 /* 0x68e0 */;
                6713: data_o = 32'h00000000 /* 0x68e4 */;
                6714: data_o = 32'h00000000 /* 0x68e8 */;
                6715: data_o = 32'h00000000 /* 0x68ec */;
                6716: data_o = 32'h00000000 /* 0x68f0 */;
                6717: data_o = 32'h00000000 /* 0x68f4 */;
                6718: data_o = 32'h00000000 /* 0x68f8 */;
                6719: data_o = 32'h00000000 /* 0x68fc */;
                6720: data_o = 32'h00000000 /* 0x6900 */;
                6721: data_o = 32'h00000000 /* 0x6904 */;
                6722: data_o = 32'h00000000 /* 0x6908 */;
                6723: data_o = 32'h00000000 /* 0x690c */;
                6724: data_o = 32'h00000000 /* 0x6910 */;
                6725: data_o = 32'h00000000 /* 0x6914 */;
                6726: data_o = 32'h00000000 /* 0x6918 */;
                6727: data_o = 32'h00000000 /* 0x691c */;
                6728: data_o = 32'h00000000 /* 0x6920 */;
                6729: data_o = 32'h00000000 /* 0x6924 */;
                6730: data_o = 32'h00000000 /* 0x6928 */;
                6731: data_o = 32'h00000000 /* 0x692c */;
                6732: data_o = 32'h00000000 /* 0x6930 */;
                6733: data_o = 32'h00000000 /* 0x6934 */;
                6734: data_o = 32'h00000000 /* 0x6938 */;
                6735: data_o = 32'h00000000 /* 0x693c */;
                6736: data_o = 32'h00000000 /* 0x6940 */;
                6737: data_o = 32'h00000000 /* 0x6944 */;
                6738: data_o = 32'h00000000 /* 0x6948 */;
                6739: data_o = 32'h00000000 /* 0x694c */;
                6740: data_o = 32'h00000000 /* 0x6950 */;
                6741: data_o = 32'h00000000 /* 0x6954 */;
                6742: data_o = 32'h00000000 /* 0x6958 */;
                6743: data_o = 32'h00000000 /* 0x695c */;
                6744: data_o = 32'h00000000 /* 0x6960 */;
                6745: data_o = 32'h00000000 /* 0x6964 */;
                6746: data_o = 32'h00000000 /* 0x6968 */;
                6747: data_o = 32'h00000000 /* 0x696c */;
                6748: data_o = 32'h00000000 /* 0x6970 */;
                6749: data_o = 32'h00000000 /* 0x6974 */;
                6750: data_o = 32'h00000000 /* 0x6978 */;
                6751: data_o = 32'h00000000 /* 0x697c */;
                6752: data_o = 32'h00000000 /* 0x6980 */;
                6753: data_o = 32'h00000000 /* 0x6984 */;
                6754: data_o = 32'h00000000 /* 0x6988 */;
                6755: data_o = 32'h00000000 /* 0x698c */;
                6756: data_o = 32'h00000000 /* 0x6990 */;
                6757: data_o = 32'h00000000 /* 0x6994 */;
                6758: data_o = 32'h00000000 /* 0x6998 */;
                6759: data_o = 32'h00000000 /* 0x699c */;
                6760: data_o = 32'h00000000 /* 0x69a0 */;
                6761: data_o = 32'h00000000 /* 0x69a4 */;
                6762: data_o = 32'h00000000 /* 0x69a8 */;
                6763: data_o = 32'h00000000 /* 0x69ac */;
                6764: data_o = 32'h00000000 /* 0x69b0 */;
                6765: data_o = 32'h00000000 /* 0x69b4 */;
                6766: data_o = 32'h00000000 /* 0x69b8 */;
                6767: data_o = 32'h00000000 /* 0x69bc */;
                6768: data_o = 32'h00000000 /* 0x69c0 */;
                6769: data_o = 32'h00000000 /* 0x69c4 */;
                6770: data_o = 32'h00000000 /* 0x69c8 */;
                6771: data_o = 32'h00000000 /* 0x69cc */;
                6772: data_o = 32'h00000000 /* 0x69d0 */;
                6773: data_o = 32'h00000000 /* 0x69d4 */;
                6774: data_o = 32'h00000000 /* 0x69d8 */;
                6775: data_o = 32'h00000000 /* 0x69dc */;
                6776: data_o = 32'h00000000 /* 0x69e0 */;
                6777: data_o = 32'h00000000 /* 0x69e4 */;
                6778: data_o = 32'h00000000 /* 0x69e8 */;
                6779: data_o = 32'h00000000 /* 0x69ec */;
                6780: data_o = 32'h00000000 /* 0x69f0 */;
                6781: data_o = 32'h00000000 /* 0x69f4 */;
                6782: data_o = 32'h00000000 /* 0x69f8 */;
                6783: data_o = 32'h00000000 /* 0x69fc */;
                6784: data_o = 32'h00000000 /* 0x6a00 */;
                6785: data_o = 32'h00000000 /* 0x6a04 */;
                6786: data_o = 32'h00000000 /* 0x6a08 */;
                6787: data_o = 32'h00000000 /* 0x6a0c */;
                6788: data_o = 32'h00000000 /* 0x6a10 */;
                6789: data_o = 32'h00000000 /* 0x6a14 */;
                6790: data_o = 32'h00000000 /* 0x6a18 */;
                6791: data_o = 32'h00000000 /* 0x6a1c */;
                6792: data_o = 32'h00000000 /* 0x6a20 */;
                6793: data_o = 32'h00000000 /* 0x6a24 */;
                6794: data_o = 32'h00000000 /* 0x6a28 */;
                6795: data_o = 32'h00000000 /* 0x6a2c */;
                6796: data_o = 32'h00000000 /* 0x6a30 */;
                6797: data_o = 32'h00000000 /* 0x6a34 */;
                6798: data_o = 32'h00000000 /* 0x6a38 */;
                6799: data_o = 32'h00000000 /* 0x6a3c */;
                6800: data_o = 32'h00000000 /* 0x6a40 */;
                6801: data_o = 32'h00000000 /* 0x6a44 */;
                6802: data_o = 32'h00000000 /* 0x6a48 */;
                6803: data_o = 32'h00000000 /* 0x6a4c */;
                6804: data_o = 32'h00000000 /* 0x6a50 */;
                6805: data_o = 32'h00000000 /* 0x6a54 */;
                6806: data_o = 32'h00000000 /* 0x6a58 */;
                6807: data_o = 32'h00000000 /* 0x6a5c */;
                6808: data_o = 32'h00000000 /* 0x6a60 */;
                6809: data_o = 32'h00000000 /* 0x6a64 */;
                6810: data_o = 32'h00000000 /* 0x6a68 */;
                6811: data_o = 32'h00000000 /* 0x6a6c */;
                6812: data_o = 32'h00000000 /* 0x6a70 */;
                6813: data_o = 32'h00000000 /* 0x6a74 */;
                6814: data_o = 32'h00000000 /* 0x6a78 */;
                6815: data_o = 32'h00000000 /* 0x6a7c */;
                6816: data_o = 32'h00000000 /* 0x6a80 */;
                6817: data_o = 32'h00000000 /* 0x6a84 */;
                6818: data_o = 32'h00000000 /* 0x6a88 */;
                6819: data_o = 32'h00000000 /* 0x6a8c */;
                6820: data_o = 32'h00000000 /* 0x6a90 */;
                6821: data_o = 32'h00000000 /* 0x6a94 */;
                6822: data_o = 32'h00000000 /* 0x6a98 */;
                6823: data_o = 32'h00000000 /* 0x6a9c */;
                6824: data_o = 32'h00000000 /* 0x6aa0 */;
                6825: data_o = 32'h00000000 /* 0x6aa4 */;
                6826: data_o = 32'h00000000 /* 0x6aa8 */;
                6827: data_o = 32'h00000000 /* 0x6aac */;
                6828: data_o = 32'h00000000 /* 0x6ab0 */;
                6829: data_o = 32'h00000000 /* 0x6ab4 */;
                6830: data_o = 32'h00000000 /* 0x6ab8 */;
                6831: data_o = 32'h00000000 /* 0x6abc */;
                6832: data_o = 32'h00000000 /* 0x6ac0 */;
                6833: data_o = 32'h00000000 /* 0x6ac4 */;
                6834: data_o = 32'h00000000 /* 0x6ac8 */;
                6835: data_o = 32'h00000000 /* 0x6acc */;
                6836: data_o = 32'h00000000 /* 0x6ad0 */;
                6837: data_o = 32'h00000000 /* 0x6ad4 */;
                6838: data_o = 32'h00000000 /* 0x6ad8 */;
                6839: data_o = 32'h00000000 /* 0x6adc */;
                6840: data_o = 32'h00000000 /* 0x6ae0 */;
                6841: data_o = 32'h00000000 /* 0x6ae4 */;
                6842: data_o = 32'h00000000 /* 0x6ae8 */;
                6843: data_o = 32'h00000000 /* 0x6aec */;
                6844: data_o = 32'h00000000 /* 0x6af0 */;
                6845: data_o = 32'h00000000 /* 0x6af4 */;
                6846: data_o = 32'h00000000 /* 0x6af8 */;
                6847: data_o = 32'h00000000 /* 0x6afc */;
                6848: data_o = 32'h00000000 /* 0x6b00 */;
                6849: data_o = 32'h00000000 /* 0x6b04 */;
                6850: data_o = 32'h00000000 /* 0x6b08 */;
                6851: data_o = 32'h00000000 /* 0x6b0c */;
                6852: data_o = 32'h00000000 /* 0x6b10 */;
                6853: data_o = 32'h00000000 /* 0x6b14 */;
                6854: data_o = 32'h00000000 /* 0x6b18 */;
                6855: data_o = 32'h00000000 /* 0x6b1c */;
                6856: data_o = 32'h00000000 /* 0x6b20 */;
                6857: data_o = 32'h00000000 /* 0x6b24 */;
                6858: data_o = 32'h00000000 /* 0x6b28 */;
                6859: data_o = 32'h00000000 /* 0x6b2c */;
                6860: data_o = 32'h00000000 /* 0x6b30 */;
                6861: data_o = 32'h00000000 /* 0x6b34 */;
                6862: data_o = 32'h00000000 /* 0x6b38 */;
                6863: data_o = 32'h00000000 /* 0x6b3c */;
                6864: data_o = 32'h00000000 /* 0x6b40 */;
                6865: data_o = 32'h00000000 /* 0x6b44 */;
                6866: data_o = 32'h00000000 /* 0x6b48 */;
                6867: data_o = 32'h00000000 /* 0x6b4c */;
                6868: data_o = 32'h00000000 /* 0x6b50 */;
                6869: data_o = 32'h00000000 /* 0x6b54 */;
                6870: data_o = 32'h00000000 /* 0x6b58 */;
                6871: data_o = 32'h00000000 /* 0x6b5c */;
                6872: data_o = 32'h00000000 /* 0x6b60 */;
                6873: data_o = 32'h00000000 /* 0x6b64 */;
                6874: data_o = 32'h00000000 /* 0x6b68 */;
                6875: data_o = 32'h00000000 /* 0x6b6c */;
                6876: data_o = 32'h00000000 /* 0x6b70 */;
                6877: data_o = 32'h00000000 /* 0x6b74 */;
                6878: data_o = 32'h00000000 /* 0x6b78 */;
                6879: data_o = 32'h00000000 /* 0x6b7c */;
                6880: data_o = 32'h00000000 /* 0x6b80 */;
                6881: data_o = 32'h00000000 /* 0x6b84 */;
                6882: data_o = 32'h00000000 /* 0x6b88 */;
                6883: data_o = 32'h00000000 /* 0x6b8c */;
                6884: data_o = 32'h00000000 /* 0x6b90 */;
                6885: data_o = 32'h00000000 /* 0x6b94 */;
                6886: data_o = 32'h00000000 /* 0x6b98 */;
                6887: data_o = 32'h00000000 /* 0x6b9c */;
                6888: data_o = 32'h00000000 /* 0x6ba0 */;
                6889: data_o = 32'h00000000 /* 0x6ba4 */;
                6890: data_o = 32'h00000000 /* 0x6ba8 */;
                6891: data_o = 32'h00000000 /* 0x6bac */;
                6892: data_o = 32'h00000000 /* 0x6bb0 */;
                6893: data_o = 32'h00000000 /* 0x6bb4 */;
                6894: data_o = 32'h00000000 /* 0x6bb8 */;
                6895: data_o = 32'h00000000 /* 0x6bbc */;
                6896: data_o = 32'h00000000 /* 0x6bc0 */;
                6897: data_o = 32'h00000000 /* 0x6bc4 */;
                6898: data_o = 32'h00000000 /* 0x6bc8 */;
                6899: data_o = 32'h00000000 /* 0x6bcc */;
                6900: data_o = 32'h00000000 /* 0x6bd0 */;
                6901: data_o = 32'h00000000 /* 0x6bd4 */;
                6902: data_o = 32'h00000000 /* 0x6bd8 */;
                6903: data_o = 32'h00000000 /* 0x6bdc */;
                6904: data_o = 32'h00000000 /* 0x6be0 */;
                6905: data_o = 32'h00000000 /* 0x6be4 */;
                6906: data_o = 32'h00000000 /* 0x6be8 */;
                6907: data_o = 32'h00000000 /* 0x6bec */;
                6908: data_o = 32'h00000000 /* 0x6bf0 */;
                6909: data_o = 32'h00000000 /* 0x6bf4 */;
                6910: data_o = 32'h00000000 /* 0x6bf8 */;
                6911: data_o = 32'h00000000 /* 0x6bfc */;
                6912: data_o = 32'h00000000 /* 0x6c00 */;
                6913: data_o = 32'h00000000 /* 0x6c04 */;
                6914: data_o = 32'h00000000 /* 0x6c08 */;
                6915: data_o = 32'h00000000 /* 0x6c0c */;
                6916: data_o = 32'h00000000 /* 0x6c10 */;
                6917: data_o = 32'h00000000 /* 0x6c14 */;
                6918: data_o = 32'h00000000 /* 0x6c18 */;
                6919: data_o = 32'h00000000 /* 0x6c1c */;
                6920: data_o = 32'h00000000 /* 0x6c20 */;
                6921: data_o = 32'h00000000 /* 0x6c24 */;
                6922: data_o = 32'h00000000 /* 0x6c28 */;
                6923: data_o = 32'h00000000 /* 0x6c2c */;
                6924: data_o = 32'h00000000 /* 0x6c30 */;
                6925: data_o = 32'h00000000 /* 0x6c34 */;
                6926: data_o = 32'h00000000 /* 0x6c38 */;
                6927: data_o = 32'h00000000 /* 0x6c3c */;
                6928: data_o = 32'h00000000 /* 0x6c40 */;
                6929: data_o = 32'h00000000 /* 0x6c44 */;
                6930: data_o = 32'h00000000 /* 0x6c48 */;
                6931: data_o = 32'h00000000 /* 0x6c4c */;
                6932: data_o = 32'h00000000 /* 0x6c50 */;
                6933: data_o = 32'h00000000 /* 0x6c54 */;
                6934: data_o = 32'h00000000 /* 0x6c58 */;
                6935: data_o = 32'h00000000 /* 0x6c5c */;
                6936: data_o = 32'h00000000 /* 0x6c60 */;
                6937: data_o = 32'h00000000 /* 0x6c64 */;
                6938: data_o = 32'h00000000 /* 0x6c68 */;
                6939: data_o = 32'h00000000 /* 0x6c6c */;
                6940: data_o = 32'h00000000 /* 0x6c70 */;
                6941: data_o = 32'h00000000 /* 0x6c74 */;
                6942: data_o = 32'h00000000 /* 0x6c78 */;
                6943: data_o = 32'h00000000 /* 0x6c7c */;
                6944: data_o = 32'h00000000 /* 0x6c80 */;
                6945: data_o = 32'h00000000 /* 0x6c84 */;
                6946: data_o = 32'h00000000 /* 0x6c88 */;
                6947: data_o = 32'h00000000 /* 0x6c8c */;
                6948: data_o = 32'h00000000 /* 0x6c90 */;
                6949: data_o = 32'h00000000 /* 0x6c94 */;
                6950: data_o = 32'h00000000 /* 0x6c98 */;
                6951: data_o = 32'h00000000 /* 0x6c9c */;
                6952: data_o = 32'h00000000 /* 0x6ca0 */;
                6953: data_o = 32'h00000000 /* 0x6ca4 */;
                6954: data_o = 32'h00000000 /* 0x6ca8 */;
                6955: data_o = 32'h00000000 /* 0x6cac */;
                6956: data_o = 32'h00000000 /* 0x6cb0 */;
                6957: data_o = 32'h00000000 /* 0x6cb4 */;
                6958: data_o = 32'h00000000 /* 0x6cb8 */;
                6959: data_o = 32'h00000000 /* 0x6cbc */;
                6960: data_o = 32'h00000000 /* 0x6cc0 */;
                6961: data_o = 32'h00000000 /* 0x6cc4 */;
                6962: data_o = 32'h00000000 /* 0x6cc8 */;
                6963: data_o = 32'h00000000 /* 0x6ccc */;
                6964: data_o = 32'h00000000 /* 0x6cd0 */;
                6965: data_o = 32'h00000000 /* 0x6cd4 */;
                6966: data_o = 32'h00000000 /* 0x6cd8 */;
                6967: data_o = 32'h00000000 /* 0x6cdc */;
                6968: data_o = 32'h00000000 /* 0x6ce0 */;
                6969: data_o = 32'h00000000 /* 0x6ce4 */;
                6970: data_o = 32'h00000000 /* 0x6ce8 */;
                6971: data_o = 32'h00000000 /* 0x6cec */;
                6972: data_o = 32'h00000000 /* 0x6cf0 */;
                6973: data_o = 32'h00000000 /* 0x6cf4 */;
                6974: data_o = 32'h00000000 /* 0x6cf8 */;
                6975: data_o = 32'h00000000 /* 0x6cfc */;
                6976: data_o = 32'h00000000 /* 0x6d00 */;
                6977: data_o = 32'h00000000 /* 0x6d04 */;
                6978: data_o = 32'h00000000 /* 0x6d08 */;
                6979: data_o = 32'h00000000 /* 0x6d0c */;
                6980: data_o = 32'h00000000 /* 0x6d10 */;
                6981: data_o = 32'h00000000 /* 0x6d14 */;
                6982: data_o = 32'h00000000 /* 0x6d18 */;
                6983: data_o = 32'h00000000 /* 0x6d1c */;
                6984: data_o = 32'h00000000 /* 0x6d20 */;
                6985: data_o = 32'h00000000 /* 0x6d24 */;
                6986: data_o = 32'h00000000 /* 0x6d28 */;
                6987: data_o = 32'h00000000 /* 0x6d2c */;
                6988: data_o = 32'h00000000 /* 0x6d30 */;
                6989: data_o = 32'h00000000 /* 0x6d34 */;
                6990: data_o = 32'h00000000 /* 0x6d38 */;
                6991: data_o = 32'h00000000 /* 0x6d3c */;
                6992: data_o = 32'h00000000 /* 0x6d40 */;
                6993: data_o = 32'h00000000 /* 0x6d44 */;
                6994: data_o = 32'h00000000 /* 0x6d48 */;
                6995: data_o = 32'h00000000 /* 0x6d4c */;
                6996: data_o = 32'h00000000 /* 0x6d50 */;
                6997: data_o = 32'h00000000 /* 0x6d54 */;
                6998: data_o = 32'h00000000 /* 0x6d58 */;
                6999: data_o = 32'h00000000 /* 0x6d5c */;
                7000: data_o = 32'h00000000 /* 0x6d60 */;
                7001: data_o = 32'h00000000 /* 0x6d64 */;
                7002: data_o = 32'h00000000 /* 0x6d68 */;
                7003: data_o = 32'h00000000 /* 0x6d6c */;
                7004: data_o = 32'h00000000 /* 0x6d70 */;
                7005: data_o = 32'h00000000 /* 0x6d74 */;
                7006: data_o = 32'h00000000 /* 0x6d78 */;
                7007: data_o = 32'h00000000 /* 0x6d7c */;
                7008: data_o = 32'h00000000 /* 0x6d80 */;
                7009: data_o = 32'h00000000 /* 0x6d84 */;
                7010: data_o = 32'h00000000 /* 0x6d88 */;
                7011: data_o = 32'h00000000 /* 0x6d8c */;
                7012: data_o = 32'h00000000 /* 0x6d90 */;
                7013: data_o = 32'h00000000 /* 0x6d94 */;
                7014: data_o = 32'h00000000 /* 0x6d98 */;
                7015: data_o = 32'h00000000 /* 0x6d9c */;
                7016: data_o = 32'h00000000 /* 0x6da0 */;
                7017: data_o = 32'h00000000 /* 0x6da4 */;
                7018: data_o = 32'h00000000 /* 0x6da8 */;
                7019: data_o = 32'h00000000 /* 0x6dac */;
                7020: data_o = 32'h00000000 /* 0x6db0 */;
                7021: data_o = 32'h00000000 /* 0x6db4 */;
                7022: data_o = 32'h00000000 /* 0x6db8 */;
                7023: data_o = 32'h00000000 /* 0x6dbc */;
                7024: data_o = 32'h00000000 /* 0x6dc0 */;
                7025: data_o = 32'h00000000 /* 0x6dc4 */;
                7026: data_o = 32'h00000000 /* 0x6dc8 */;
                7027: data_o = 32'h00000000 /* 0x6dcc */;
                7028: data_o = 32'h00000000 /* 0x6dd0 */;
                7029: data_o = 32'h00000000 /* 0x6dd4 */;
                7030: data_o = 32'h00000000 /* 0x6dd8 */;
                7031: data_o = 32'h00000000 /* 0x6ddc */;
                7032: data_o = 32'h00000000 /* 0x6de0 */;
                7033: data_o = 32'h00000000 /* 0x6de4 */;
                7034: data_o = 32'h00000000 /* 0x6de8 */;
                7035: data_o = 32'h00000000 /* 0x6dec */;
                7036: data_o = 32'h00000000 /* 0x6df0 */;
                7037: data_o = 32'h00000000 /* 0x6df4 */;
                7038: data_o = 32'h00000000 /* 0x6df8 */;
                7039: data_o = 32'h00000000 /* 0x6dfc */;
                7040: data_o = 32'h00000000 /* 0x6e00 */;
                7041: data_o = 32'h00000000 /* 0x6e04 */;
                7042: data_o = 32'h00000000 /* 0x6e08 */;
                7043: data_o = 32'h00000000 /* 0x6e0c */;
                7044: data_o = 32'h00000000 /* 0x6e10 */;
                7045: data_o = 32'h00000000 /* 0x6e14 */;
                7046: data_o = 32'h00000000 /* 0x6e18 */;
                7047: data_o = 32'h00000000 /* 0x6e1c */;
                7048: data_o = 32'h00000000 /* 0x6e20 */;
                7049: data_o = 32'h00000000 /* 0x6e24 */;
                7050: data_o = 32'h00000000 /* 0x6e28 */;
                7051: data_o = 32'h00000000 /* 0x6e2c */;
                7052: data_o = 32'h00000000 /* 0x6e30 */;
                7053: data_o = 32'h00000000 /* 0x6e34 */;
                7054: data_o = 32'h00000000 /* 0x6e38 */;
                7055: data_o = 32'h00000000 /* 0x6e3c */;
                7056: data_o = 32'h00000000 /* 0x6e40 */;
                7057: data_o = 32'h00000000 /* 0x6e44 */;
                7058: data_o = 32'h00000000 /* 0x6e48 */;
                7059: data_o = 32'h00000000 /* 0x6e4c */;
                7060: data_o = 32'h00000000 /* 0x6e50 */;
                7061: data_o = 32'h00000000 /* 0x6e54 */;
                7062: data_o = 32'h00000000 /* 0x6e58 */;
                7063: data_o = 32'h00000000 /* 0x6e5c */;
                7064: data_o = 32'h00000000 /* 0x6e60 */;
                7065: data_o = 32'h00000000 /* 0x6e64 */;
                7066: data_o = 32'h00000000 /* 0x6e68 */;
                7067: data_o = 32'h00000000 /* 0x6e6c */;
                7068: data_o = 32'h00000000 /* 0x6e70 */;
                7069: data_o = 32'h00000000 /* 0x6e74 */;
                7070: data_o = 32'h00000000 /* 0x6e78 */;
                7071: data_o = 32'h00000000 /* 0x6e7c */;
                7072: data_o = 32'h00000000 /* 0x6e80 */;
                7073: data_o = 32'h00000000 /* 0x6e84 */;
                7074: data_o = 32'h00000000 /* 0x6e88 */;
                7075: data_o = 32'h00000000 /* 0x6e8c */;
                7076: data_o = 32'h00000000 /* 0x6e90 */;
                7077: data_o = 32'h00000000 /* 0x6e94 */;
                7078: data_o = 32'h00000000 /* 0x6e98 */;
                7079: data_o = 32'h00000000 /* 0x6e9c */;
                7080: data_o = 32'h00000000 /* 0x6ea0 */;
                7081: data_o = 32'h00000000 /* 0x6ea4 */;
                7082: data_o = 32'h00000000 /* 0x6ea8 */;
                7083: data_o = 32'h00000000 /* 0x6eac */;
                7084: data_o = 32'h00000000 /* 0x6eb0 */;
                7085: data_o = 32'h00000000 /* 0x6eb4 */;
                7086: data_o = 32'h00000000 /* 0x6eb8 */;
                7087: data_o = 32'h00000000 /* 0x6ebc */;
                7088: data_o = 32'h00000000 /* 0x6ec0 */;
                7089: data_o = 32'h00000000 /* 0x6ec4 */;
                7090: data_o = 32'h00000000 /* 0x6ec8 */;
                7091: data_o = 32'h00000000 /* 0x6ecc */;
                7092: data_o = 32'h00000000 /* 0x6ed0 */;
                7093: data_o = 32'h00000000 /* 0x6ed4 */;
                7094: data_o = 32'h00000000 /* 0x6ed8 */;
                7095: data_o = 32'h00000000 /* 0x6edc */;
                7096: data_o = 32'h00000000 /* 0x6ee0 */;
                7097: data_o = 32'h00000000 /* 0x6ee4 */;
                7098: data_o = 32'h00000000 /* 0x6ee8 */;
                7099: data_o = 32'h00000000 /* 0x6eec */;
                7100: data_o = 32'h00000000 /* 0x6ef0 */;
                7101: data_o = 32'h00000000 /* 0x6ef4 */;
                7102: data_o = 32'h00000000 /* 0x6ef8 */;
                7103: data_o = 32'h00000000 /* 0x6efc */;
                7104: data_o = 32'h00000000 /* 0x6f00 */;
                7105: data_o = 32'h00000000 /* 0x6f04 */;
                7106: data_o = 32'h00000000 /* 0x6f08 */;
                7107: data_o = 32'h00000000 /* 0x6f0c */;
                7108: data_o = 32'h00000000 /* 0x6f10 */;
                7109: data_o = 32'h00000000 /* 0x6f14 */;
                7110: data_o = 32'h00000000 /* 0x6f18 */;
                7111: data_o = 32'h00000000 /* 0x6f1c */;
                7112: data_o = 32'h00000000 /* 0x6f20 */;
                7113: data_o = 32'h00000000 /* 0x6f24 */;
                7114: data_o = 32'h00000000 /* 0x6f28 */;
                7115: data_o = 32'h00000000 /* 0x6f2c */;
                7116: data_o = 32'h00000000 /* 0x6f30 */;
                7117: data_o = 32'h00000000 /* 0x6f34 */;
                7118: data_o = 32'h00000000 /* 0x6f38 */;
                7119: data_o = 32'h00000000 /* 0x6f3c */;
                7120: data_o = 32'h00000000 /* 0x6f40 */;
                7121: data_o = 32'h00000000 /* 0x6f44 */;
                7122: data_o = 32'h00000000 /* 0x6f48 */;
                7123: data_o = 32'h00000000 /* 0x6f4c */;
                7124: data_o = 32'h00000000 /* 0x6f50 */;
                7125: data_o = 32'h00000000 /* 0x6f54 */;
                7126: data_o = 32'h00000000 /* 0x6f58 */;
                7127: data_o = 32'h00000000 /* 0x6f5c */;
                7128: data_o = 32'h00000000 /* 0x6f60 */;
                7129: data_o = 32'h00000000 /* 0x6f64 */;
                7130: data_o = 32'h00000000 /* 0x6f68 */;
                7131: data_o = 32'h00000000 /* 0x6f6c */;
                7132: data_o = 32'h00000000 /* 0x6f70 */;
                7133: data_o = 32'h00000000 /* 0x6f74 */;
                7134: data_o = 32'h00000000 /* 0x6f78 */;
                7135: data_o = 32'h00000000 /* 0x6f7c */;
                7136: data_o = 32'h00000000 /* 0x6f80 */;
                7137: data_o = 32'h00000000 /* 0x6f84 */;
                7138: data_o = 32'h00000000 /* 0x6f88 */;
                7139: data_o = 32'h00000000 /* 0x6f8c */;
                7140: data_o = 32'h00000000 /* 0x6f90 */;
                7141: data_o = 32'h00000000 /* 0x6f94 */;
                7142: data_o = 32'h00000000 /* 0x6f98 */;
                7143: data_o = 32'h00000000 /* 0x6f9c */;
                7144: data_o = 32'h00000000 /* 0x6fa0 */;
                7145: data_o = 32'h00000000 /* 0x6fa4 */;
                7146: data_o = 32'h00000000 /* 0x6fa8 */;
                7147: data_o = 32'h00000000 /* 0x6fac */;
                7148: data_o = 32'h00000000 /* 0x6fb0 */;
                7149: data_o = 32'h00000000 /* 0x6fb4 */;
                7150: data_o = 32'h00000000 /* 0x6fb8 */;
                7151: data_o = 32'h00000000 /* 0x6fbc */;
                7152: data_o = 32'h00000000 /* 0x6fc0 */;
                7153: data_o = 32'h00000000 /* 0x6fc4 */;
                7154: data_o = 32'h00000000 /* 0x6fc8 */;
                7155: data_o = 32'h00000000 /* 0x6fcc */;
                7156: data_o = 32'h00000000 /* 0x6fd0 */;
                7157: data_o = 32'h00000000 /* 0x6fd4 */;
                7158: data_o = 32'h00000000 /* 0x6fd8 */;
                7159: data_o = 32'h00000000 /* 0x6fdc */;
                7160: data_o = 32'h00000000 /* 0x6fe0 */;
                7161: data_o = 32'h00000000 /* 0x6fe4 */;
                7162: data_o = 32'h00000000 /* 0x6fe8 */;
                7163: data_o = 32'h00000000 /* 0x6fec */;
                7164: data_o = 32'h00000000 /* 0x6ff0 */;
                7165: data_o = 32'h00000000 /* 0x6ff4 */;
                7166: data_o = 32'h00000000 /* 0x6ff8 */;
                7167: data_o = 32'h00000000 /* 0x6ffc */;
                7168: data_o = 32'h00000000 /* 0x7000 */;
                7169: data_o = 32'h00000000 /* 0x7004 */;
                7170: data_o = 32'h00000000 /* 0x7008 */;
                7171: data_o = 32'h00000000 /* 0x700c */;
                7172: data_o = 32'h00000000 /* 0x7010 */;
                7173: data_o = 32'h00000000 /* 0x7014 */;
                7174: data_o = 32'h00000000 /* 0x7018 */;
                7175: data_o = 32'h00000000 /* 0x701c */;
                7176: data_o = 32'h00000000 /* 0x7020 */;
                7177: data_o = 32'h00000000 /* 0x7024 */;
                7178: data_o = 32'h00000000 /* 0x7028 */;
                7179: data_o = 32'h00000000 /* 0x702c */;
                7180: data_o = 32'h00000000 /* 0x7030 */;
                7181: data_o = 32'h00000000 /* 0x7034 */;
                7182: data_o = 32'h00000000 /* 0x7038 */;
                7183: data_o = 32'h00000000 /* 0x703c */;
                7184: data_o = 32'h00000000 /* 0x7040 */;
                7185: data_o = 32'h00000000 /* 0x7044 */;
                7186: data_o = 32'h00000000 /* 0x7048 */;
                7187: data_o = 32'h00000000 /* 0x704c */;
                7188: data_o = 32'h00000000 /* 0x7050 */;
                7189: data_o = 32'h00000000 /* 0x7054 */;
                7190: data_o = 32'h00000000 /* 0x7058 */;
                7191: data_o = 32'h00000000 /* 0x705c */;
                7192: data_o = 32'h00000000 /* 0x7060 */;
                7193: data_o = 32'h00000000 /* 0x7064 */;
                7194: data_o = 32'h00000000 /* 0x7068 */;
                7195: data_o = 32'h00000000 /* 0x706c */;
                7196: data_o = 32'h00000000 /* 0x7070 */;
                7197: data_o = 32'h00000000 /* 0x7074 */;
                7198: data_o = 32'h00000000 /* 0x7078 */;
                7199: data_o = 32'h00000000 /* 0x707c */;
                7200: data_o = 32'h00000000 /* 0x7080 */;
                7201: data_o = 32'h00000000 /* 0x7084 */;
                7202: data_o = 32'h00000000 /* 0x7088 */;
                7203: data_o = 32'h00000000 /* 0x708c */;
                7204: data_o = 32'h00000000 /* 0x7090 */;
                7205: data_o = 32'h00000000 /* 0x7094 */;
                7206: data_o = 32'h00000000 /* 0x7098 */;
                7207: data_o = 32'h00000000 /* 0x709c */;
                7208: data_o = 32'h00000000 /* 0x70a0 */;
                7209: data_o = 32'h00000000 /* 0x70a4 */;
                7210: data_o = 32'h00000000 /* 0x70a8 */;
                7211: data_o = 32'h00000000 /* 0x70ac */;
                7212: data_o = 32'h00000000 /* 0x70b0 */;
                7213: data_o = 32'h00000000 /* 0x70b4 */;
                7214: data_o = 32'h00000000 /* 0x70b8 */;
                7215: data_o = 32'h00000000 /* 0x70bc */;
                7216: data_o = 32'h00000000 /* 0x70c0 */;
                7217: data_o = 32'h00000000 /* 0x70c4 */;
                7218: data_o = 32'h00000000 /* 0x70c8 */;
                7219: data_o = 32'h00000000 /* 0x70cc */;
                7220: data_o = 32'h00000000 /* 0x70d0 */;
                7221: data_o = 32'h00000000 /* 0x70d4 */;
                7222: data_o = 32'h00000000 /* 0x70d8 */;
                7223: data_o = 32'h00000000 /* 0x70dc */;
                7224: data_o = 32'h00000000 /* 0x70e0 */;
                7225: data_o = 32'h00000000 /* 0x70e4 */;
                7226: data_o = 32'h00000000 /* 0x70e8 */;
                7227: data_o = 32'h00000000 /* 0x70ec */;
                7228: data_o = 32'h00000000 /* 0x70f0 */;
                7229: data_o = 32'h00000000 /* 0x70f4 */;
                7230: data_o = 32'h00000000 /* 0x70f8 */;
                7231: data_o = 32'h00000000 /* 0x70fc */;
                7232: data_o = 32'h00000000 /* 0x7100 */;
                7233: data_o = 32'h00000000 /* 0x7104 */;
                7234: data_o = 32'h00000000 /* 0x7108 */;
                7235: data_o = 32'h00000000 /* 0x710c */;
                7236: data_o = 32'h00000000 /* 0x7110 */;
                7237: data_o = 32'h00000000 /* 0x7114 */;
                7238: data_o = 32'h00000000 /* 0x7118 */;
                7239: data_o = 32'h00000000 /* 0x711c */;
                7240: data_o = 32'h00000000 /* 0x7120 */;
                7241: data_o = 32'h00000000 /* 0x7124 */;
                7242: data_o = 32'h00000000 /* 0x7128 */;
                7243: data_o = 32'h00000000 /* 0x712c */;
                7244: data_o = 32'h00000000 /* 0x7130 */;
                7245: data_o = 32'h00000000 /* 0x7134 */;
                7246: data_o = 32'h00000000 /* 0x7138 */;
                7247: data_o = 32'h00000000 /* 0x713c */;
                7248: data_o = 32'h00000000 /* 0x7140 */;
                7249: data_o = 32'h00000000 /* 0x7144 */;
                7250: data_o = 32'h00000000 /* 0x7148 */;
                7251: data_o = 32'h00000000 /* 0x714c */;
                7252: data_o = 32'h00000000 /* 0x7150 */;
                7253: data_o = 32'h00000000 /* 0x7154 */;
                7254: data_o = 32'h00000000 /* 0x7158 */;
                7255: data_o = 32'h00000000 /* 0x715c */;
                7256: data_o = 32'h00000000 /* 0x7160 */;
                7257: data_o = 32'h00000000 /* 0x7164 */;
                7258: data_o = 32'h00000000 /* 0x7168 */;
                7259: data_o = 32'h00000000 /* 0x716c */;
                7260: data_o = 32'h00000000 /* 0x7170 */;
                7261: data_o = 32'h00000000 /* 0x7174 */;
                7262: data_o = 32'h00000000 /* 0x7178 */;
                7263: data_o = 32'h00000000 /* 0x717c */;
                7264: data_o = 32'h00000000 /* 0x7180 */;
                7265: data_o = 32'h00000000 /* 0x7184 */;
                7266: data_o = 32'h00000000 /* 0x7188 */;
                7267: data_o = 32'h00000000 /* 0x718c */;
                7268: data_o = 32'h00000000 /* 0x7190 */;
                7269: data_o = 32'h00000000 /* 0x7194 */;
                7270: data_o = 32'h00000000 /* 0x7198 */;
                7271: data_o = 32'h00000000 /* 0x719c */;
                7272: data_o = 32'h00000000 /* 0x71a0 */;
                7273: data_o = 32'h00000000 /* 0x71a4 */;
                7274: data_o = 32'h00000000 /* 0x71a8 */;
                7275: data_o = 32'h00000000 /* 0x71ac */;
                7276: data_o = 32'h00000000 /* 0x71b0 */;
                7277: data_o = 32'h00000000 /* 0x71b4 */;
                7278: data_o = 32'h00000000 /* 0x71b8 */;
                7279: data_o = 32'h00000000 /* 0x71bc */;
                7280: data_o = 32'h00000000 /* 0x71c0 */;
                7281: data_o = 32'h00000000 /* 0x71c4 */;
                7282: data_o = 32'h00000000 /* 0x71c8 */;
                7283: data_o = 32'h00000000 /* 0x71cc */;
                7284: data_o = 32'h00000000 /* 0x71d0 */;
                7285: data_o = 32'h00000000 /* 0x71d4 */;
                7286: data_o = 32'h00000000 /* 0x71d8 */;
                7287: data_o = 32'h00000000 /* 0x71dc */;
                7288: data_o = 32'h00000000 /* 0x71e0 */;
                7289: data_o = 32'h00000000 /* 0x71e4 */;
                7290: data_o = 32'h00000000 /* 0x71e8 */;
                7291: data_o = 32'h00000000 /* 0x71ec */;
                7292: data_o = 32'h00000000 /* 0x71f0 */;
                7293: data_o = 32'h00000000 /* 0x71f4 */;
                7294: data_o = 32'h00000000 /* 0x71f8 */;
                7295: data_o = 32'h00000000 /* 0x71fc */;
                7296: data_o = 32'h00000000 /* 0x7200 */;
                7297: data_o = 32'h00000000 /* 0x7204 */;
                7298: data_o = 32'h00000000 /* 0x7208 */;
                7299: data_o = 32'h00000000 /* 0x720c */;
                7300: data_o = 32'h00000000 /* 0x7210 */;
                7301: data_o = 32'h00000000 /* 0x7214 */;
                7302: data_o = 32'h00000000 /* 0x7218 */;
                7303: data_o = 32'h00000000 /* 0x721c */;
                7304: data_o = 32'h00000000 /* 0x7220 */;
                7305: data_o = 32'h00000000 /* 0x7224 */;
                7306: data_o = 32'h00000000 /* 0x7228 */;
                7307: data_o = 32'h00000000 /* 0x722c */;
                7308: data_o = 32'h00000000 /* 0x7230 */;
                7309: data_o = 32'h00000000 /* 0x7234 */;
                7310: data_o = 32'h00000000 /* 0x7238 */;
                7311: data_o = 32'h00000000 /* 0x723c */;
                7312: data_o = 32'h00000000 /* 0x7240 */;
                7313: data_o = 32'h00000000 /* 0x7244 */;
                7314: data_o = 32'h00000000 /* 0x7248 */;
                7315: data_o = 32'h00000000 /* 0x724c */;
                7316: data_o = 32'h00000000 /* 0x7250 */;
                7317: data_o = 32'h00000000 /* 0x7254 */;
                7318: data_o = 32'h00000000 /* 0x7258 */;
                7319: data_o = 32'h00000000 /* 0x725c */;
                7320: data_o = 32'h00000000 /* 0x7260 */;
                7321: data_o = 32'h00000000 /* 0x7264 */;
                7322: data_o = 32'h00000000 /* 0x7268 */;
                7323: data_o = 32'h00000000 /* 0x726c */;
                7324: data_o = 32'h00000000 /* 0x7270 */;
                7325: data_o = 32'h00000000 /* 0x7274 */;
                7326: data_o = 32'h00000000 /* 0x7278 */;
                7327: data_o = 32'h00000000 /* 0x727c */;
                7328: data_o = 32'h00000000 /* 0x7280 */;
                7329: data_o = 32'h00000000 /* 0x7284 */;
                7330: data_o = 32'h00000000 /* 0x7288 */;
                7331: data_o = 32'h00000000 /* 0x728c */;
                7332: data_o = 32'h00000000 /* 0x7290 */;
                7333: data_o = 32'h00000000 /* 0x7294 */;
                7334: data_o = 32'h00000000 /* 0x7298 */;
                7335: data_o = 32'h00000000 /* 0x729c */;
                7336: data_o = 32'h00000000 /* 0x72a0 */;
                7337: data_o = 32'h00000000 /* 0x72a4 */;
                7338: data_o = 32'h00000000 /* 0x72a8 */;
                7339: data_o = 32'h00000000 /* 0x72ac */;
                7340: data_o = 32'h00000000 /* 0x72b0 */;
                7341: data_o = 32'h00000000 /* 0x72b4 */;
                7342: data_o = 32'h00000000 /* 0x72b8 */;
                7343: data_o = 32'h00000000 /* 0x72bc */;
                7344: data_o = 32'h00000000 /* 0x72c0 */;
                7345: data_o = 32'h00000000 /* 0x72c4 */;
                7346: data_o = 32'h00000000 /* 0x72c8 */;
                7347: data_o = 32'h00000000 /* 0x72cc */;
                7348: data_o = 32'h00000000 /* 0x72d0 */;
                7349: data_o = 32'h00000000 /* 0x72d4 */;
                7350: data_o = 32'h00000000 /* 0x72d8 */;
                7351: data_o = 32'h00000000 /* 0x72dc */;
                7352: data_o = 32'h00000000 /* 0x72e0 */;
                7353: data_o = 32'h00000000 /* 0x72e4 */;
                7354: data_o = 32'h00000000 /* 0x72e8 */;
                7355: data_o = 32'h00000000 /* 0x72ec */;
                7356: data_o = 32'h00000000 /* 0x72f0 */;
                7357: data_o = 32'h00000000 /* 0x72f4 */;
                7358: data_o = 32'h00000000 /* 0x72f8 */;
                7359: data_o = 32'h00000000 /* 0x72fc */;
                7360: data_o = 32'h00000000 /* 0x7300 */;
                7361: data_o = 32'h00000000 /* 0x7304 */;
                7362: data_o = 32'h00000000 /* 0x7308 */;
                7363: data_o = 32'h00000000 /* 0x730c */;
                7364: data_o = 32'h00000000 /* 0x7310 */;
                7365: data_o = 32'h00000000 /* 0x7314 */;
                7366: data_o = 32'h00000000 /* 0x7318 */;
                7367: data_o = 32'h00000000 /* 0x731c */;
                7368: data_o = 32'h00000000 /* 0x7320 */;
                7369: data_o = 32'h00000000 /* 0x7324 */;
                7370: data_o = 32'h00000000 /* 0x7328 */;
                7371: data_o = 32'h00000000 /* 0x732c */;
                7372: data_o = 32'h00000000 /* 0x7330 */;
                7373: data_o = 32'h00000000 /* 0x7334 */;
                7374: data_o = 32'h00000000 /* 0x7338 */;
                7375: data_o = 32'h00000000 /* 0x733c */;
                7376: data_o = 32'h00000000 /* 0x7340 */;
                7377: data_o = 32'h00000000 /* 0x7344 */;
                7378: data_o = 32'h00000000 /* 0x7348 */;
                7379: data_o = 32'h00000000 /* 0x734c */;
                7380: data_o = 32'h00000000 /* 0x7350 */;
                7381: data_o = 32'h00000000 /* 0x7354 */;
                7382: data_o = 32'h00000000 /* 0x7358 */;
                7383: data_o = 32'h00000000 /* 0x735c */;
                7384: data_o = 32'h00000000 /* 0x7360 */;
                7385: data_o = 32'h00000000 /* 0x7364 */;
                7386: data_o = 32'h00000000 /* 0x7368 */;
                7387: data_o = 32'h00000000 /* 0x736c */;
                7388: data_o = 32'h00000000 /* 0x7370 */;
                7389: data_o = 32'h00000000 /* 0x7374 */;
                7390: data_o = 32'h00000000 /* 0x7378 */;
                7391: data_o = 32'h00000000 /* 0x737c */;
                7392: data_o = 32'h00000000 /* 0x7380 */;
                7393: data_o = 32'h00000000 /* 0x7384 */;
                7394: data_o = 32'h00000000 /* 0x7388 */;
                7395: data_o = 32'h00000000 /* 0x738c */;
                7396: data_o = 32'h00000000 /* 0x7390 */;
                7397: data_o = 32'h00000000 /* 0x7394 */;
                7398: data_o = 32'h00000000 /* 0x7398 */;
                7399: data_o = 32'h00000000 /* 0x739c */;
                7400: data_o = 32'h00000000 /* 0x73a0 */;
                7401: data_o = 32'h00000000 /* 0x73a4 */;
                7402: data_o = 32'h00000000 /* 0x73a8 */;
                7403: data_o = 32'h00000000 /* 0x73ac */;
                7404: data_o = 32'h00000000 /* 0x73b0 */;
                7405: data_o = 32'h00000000 /* 0x73b4 */;
                7406: data_o = 32'h00000000 /* 0x73b8 */;
                7407: data_o = 32'h00000000 /* 0x73bc */;
                7408: data_o = 32'h00000000 /* 0x73c0 */;
                7409: data_o = 32'h00000000 /* 0x73c4 */;
                7410: data_o = 32'h00000000 /* 0x73c8 */;
                7411: data_o = 32'h00000000 /* 0x73cc */;
                7412: data_o = 32'h00000000 /* 0x73d0 */;
                7413: data_o = 32'h00000000 /* 0x73d4 */;
                7414: data_o = 32'h00000000 /* 0x73d8 */;
                7415: data_o = 32'h00000000 /* 0x73dc */;
                7416: data_o = 32'h00000000 /* 0x73e0 */;
                7417: data_o = 32'h00000000 /* 0x73e4 */;
                7418: data_o = 32'h00000000 /* 0x73e8 */;
                7419: data_o = 32'h00000000 /* 0x73ec */;
                7420: data_o = 32'h00000000 /* 0x73f0 */;
                7421: data_o = 32'h00000000 /* 0x73f4 */;
                7422: data_o = 32'h00000000 /* 0x73f8 */;
                7423: data_o = 32'h00000000 /* 0x73fc */;
                7424: data_o = 32'h00000000 /* 0x7400 */;
                7425: data_o = 32'h00000000 /* 0x7404 */;
                7426: data_o = 32'h00000000 /* 0x7408 */;
                7427: data_o = 32'h00000000 /* 0x740c */;
                7428: data_o = 32'h00000000 /* 0x7410 */;
                7429: data_o = 32'h00000000 /* 0x7414 */;
                7430: data_o = 32'h00000000 /* 0x7418 */;
                7431: data_o = 32'h00000000 /* 0x741c */;
                7432: data_o = 32'h00000000 /* 0x7420 */;
                7433: data_o = 32'h00000000 /* 0x7424 */;
                7434: data_o = 32'h00000000 /* 0x7428 */;
                7435: data_o = 32'h00000000 /* 0x742c */;
                7436: data_o = 32'h00000000 /* 0x7430 */;
                7437: data_o = 32'h00000000 /* 0x7434 */;
                7438: data_o = 32'h00000000 /* 0x7438 */;
                7439: data_o = 32'h00000000 /* 0x743c */;
                7440: data_o = 32'h00000000 /* 0x7440 */;
                7441: data_o = 32'h00000000 /* 0x7444 */;
                7442: data_o = 32'h00000000 /* 0x7448 */;
                7443: data_o = 32'h00000000 /* 0x744c */;
                7444: data_o = 32'h00000000 /* 0x7450 */;
                7445: data_o = 32'h00000000 /* 0x7454 */;
                7446: data_o = 32'h00000000 /* 0x7458 */;
                7447: data_o = 32'h00000000 /* 0x745c */;
                7448: data_o = 32'h00000000 /* 0x7460 */;
                7449: data_o = 32'h00000000 /* 0x7464 */;
                7450: data_o = 32'h00000000 /* 0x7468 */;
                7451: data_o = 32'h00000000 /* 0x746c */;
                7452: data_o = 32'h00000000 /* 0x7470 */;
                7453: data_o = 32'h00000000 /* 0x7474 */;
                7454: data_o = 32'h00000000 /* 0x7478 */;
                7455: data_o = 32'h00000000 /* 0x747c */;
                7456: data_o = 32'h00000000 /* 0x7480 */;
                7457: data_o = 32'h00000000 /* 0x7484 */;
                7458: data_o = 32'h00000000 /* 0x7488 */;
                7459: data_o = 32'h00000000 /* 0x748c */;
                7460: data_o = 32'h00000000 /* 0x7490 */;
                7461: data_o = 32'h00000000 /* 0x7494 */;
                7462: data_o = 32'h00000000 /* 0x7498 */;
                7463: data_o = 32'h00000000 /* 0x749c */;
                7464: data_o = 32'h00000000 /* 0x74a0 */;
                7465: data_o = 32'h00000000 /* 0x74a4 */;
                7466: data_o = 32'h00000000 /* 0x74a8 */;
                7467: data_o = 32'h00000000 /* 0x74ac */;
                7468: data_o = 32'h00000000 /* 0x74b0 */;
                7469: data_o = 32'h00000000 /* 0x74b4 */;
                7470: data_o = 32'h00000000 /* 0x74b8 */;
                7471: data_o = 32'h00000000 /* 0x74bc */;
                7472: data_o = 32'h00000000 /* 0x74c0 */;
                7473: data_o = 32'h00000000 /* 0x74c4 */;
                7474: data_o = 32'h00000000 /* 0x74c8 */;
                7475: data_o = 32'h00000000 /* 0x74cc */;
                7476: data_o = 32'h00000000 /* 0x74d0 */;
                7477: data_o = 32'h00000000 /* 0x74d4 */;
                7478: data_o = 32'h00000000 /* 0x74d8 */;
                7479: data_o = 32'h00000000 /* 0x74dc */;
                7480: data_o = 32'h00000000 /* 0x74e0 */;
                7481: data_o = 32'h00000000 /* 0x74e4 */;
                7482: data_o = 32'h00000000 /* 0x74e8 */;
                7483: data_o = 32'h00000000 /* 0x74ec */;
                7484: data_o = 32'h00000000 /* 0x74f0 */;
                7485: data_o = 32'h00000000 /* 0x74f4 */;
                7486: data_o = 32'h00000000 /* 0x74f8 */;
                7487: data_o = 32'h00000000 /* 0x74fc */;
                7488: data_o = 32'h00000000 /* 0x7500 */;
                7489: data_o = 32'h00000000 /* 0x7504 */;
                7490: data_o = 32'h00000000 /* 0x7508 */;
                7491: data_o = 32'h00000000 /* 0x750c */;
                7492: data_o = 32'h00000000 /* 0x7510 */;
                7493: data_o = 32'h00000000 /* 0x7514 */;
                7494: data_o = 32'h00000000 /* 0x7518 */;
                7495: data_o = 32'h00000000 /* 0x751c */;
                7496: data_o = 32'h00000000 /* 0x7520 */;
                7497: data_o = 32'h00000000 /* 0x7524 */;
                7498: data_o = 32'h00000000 /* 0x7528 */;
                7499: data_o = 32'h00000000 /* 0x752c */;
                7500: data_o = 32'h00000000 /* 0x7530 */;
                7501: data_o = 32'h00000000 /* 0x7534 */;
                7502: data_o = 32'h00000000 /* 0x7538 */;
                7503: data_o = 32'h00000000 /* 0x753c */;
                7504: data_o = 32'h00000000 /* 0x7540 */;
                7505: data_o = 32'h00000000 /* 0x7544 */;
                7506: data_o = 32'h00000000 /* 0x7548 */;
                7507: data_o = 32'h00000000 /* 0x754c */;
                7508: data_o = 32'h00000000 /* 0x7550 */;
                7509: data_o = 32'h00000000 /* 0x7554 */;
                7510: data_o = 32'h00000000 /* 0x7558 */;
                7511: data_o = 32'h00000000 /* 0x755c */;
                7512: data_o = 32'h00000000 /* 0x7560 */;
                7513: data_o = 32'h00000000 /* 0x7564 */;
                7514: data_o = 32'h00000000 /* 0x7568 */;
                7515: data_o = 32'h00000000 /* 0x756c */;
                7516: data_o = 32'h00000000 /* 0x7570 */;
                7517: data_o = 32'h00000000 /* 0x7574 */;
                7518: data_o = 32'h00000000 /* 0x7578 */;
                7519: data_o = 32'h00000000 /* 0x757c */;
                7520: data_o = 32'h00000000 /* 0x7580 */;
                7521: data_o = 32'h00000000 /* 0x7584 */;
                7522: data_o = 32'h00000000 /* 0x7588 */;
                7523: data_o = 32'h00000000 /* 0x758c */;
                7524: data_o = 32'h00000000 /* 0x7590 */;
                7525: data_o = 32'h00000000 /* 0x7594 */;
                7526: data_o = 32'h00000000 /* 0x7598 */;
                7527: data_o = 32'h00000000 /* 0x759c */;
                7528: data_o = 32'h00000000 /* 0x75a0 */;
                7529: data_o = 32'h00000000 /* 0x75a4 */;
                7530: data_o = 32'h00000000 /* 0x75a8 */;
                7531: data_o = 32'h00000000 /* 0x75ac */;
                7532: data_o = 32'h00000000 /* 0x75b0 */;
                7533: data_o = 32'h00000000 /* 0x75b4 */;
                7534: data_o = 32'h00000000 /* 0x75b8 */;
                7535: data_o = 32'h00000000 /* 0x75bc */;
                7536: data_o = 32'h00000000 /* 0x75c0 */;
                7537: data_o = 32'h00000000 /* 0x75c4 */;
                7538: data_o = 32'h00000000 /* 0x75c8 */;
                7539: data_o = 32'h00000000 /* 0x75cc */;
                7540: data_o = 32'h00000000 /* 0x75d0 */;
                7541: data_o = 32'h00000000 /* 0x75d4 */;
                7542: data_o = 32'h00000000 /* 0x75d8 */;
                7543: data_o = 32'h00000000 /* 0x75dc */;
                7544: data_o = 32'h00000000 /* 0x75e0 */;
                7545: data_o = 32'h00000000 /* 0x75e4 */;
                7546: data_o = 32'h00000000 /* 0x75e8 */;
                7547: data_o = 32'h00000000 /* 0x75ec */;
                7548: data_o = 32'h00000000 /* 0x75f0 */;
                7549: data_o = 32'h00000000 /* 0x75f4 */;
                7550: data_o = 32'h00000000 /* 0x75f8 */;
                7551: data_o = 32'h00000000 /* 0x75fc */;
                7552: data_o = 32'h00000000 /* 0x7600 */;
                7553: data_o = 32'h00000000 /* 0x7604 */;
                7554: data_o = 32'h00000000 /* 0x7608 */;
                7555: data_o = 32'h00000000 /* 0x760c */;
                7556: data_o = 32'h00000000 /* 0x7610 */;
                7557: data_o = 32'h00000000 /* 0x7614 */;
                7558: data_o = 32'h00000000 /* 0x7618 */;
                7559: data_o = 32'h00000000 /* 0x761c */;
                7560: data_o = 32'h00000000 /* 0x7620 */;
                7561: data_o = 32'h00000000 /* 0x7624 */;
                7562: data_o = 32'h00000000 /* 0x7628 */;
                7563: data_o = 32'h00000000 /* 0x762c */;
                7564: data_o = 32'h00000000 /* 0x7630 */;
                7565: data_o = 32'h00000000 /* 0x7634 */;
                7566: data_o = 32'h00000000 /* 0x7638 */;
                7567: data_o = 32'h00000000 /* 0x763c */;
                7568: data_o = 32'h00000000 /* 0x7640 */;
                7569: data_o = 32'h00000000 /* 0x7644 */;
                7570: data_o = 32'h00000000 /* 0x7648 */;
                7571: data_o = 32'h00000000 /* 0x764c */;
                7572: data_o = 32'h00000000 /* 0x7650 */;
                7573: data_o = 32'h00000000 /* 0x7654 */;
                7574: data_o = 32'h00000000 /* 0x7658 */;
                7575: data_o = 32'h00000000 /* 0x765c */;
                7576: data_o = 32'h00000000 /* 0x7660 */;
                7577: data_o = 32'h00000000 /* 0x7664 */;
                7578: data_o = 32'h00000000 /* 0x7668 */;
                7579: data_o = 32'h00000000 /* 0x766c */;
                7580: data_o = 32'h00000000 /* 0x7670 */;
                7581: data_o = 32'h00000000 /* 0x7674 */;
                7582: data_o = 32'h00000000 /* 0x7678 */;
                7583: data_o = 32'h00000000 /* 0x767c */;
                7584: data_o = 32'h00000000 /* 0x7680 */;
                7585: data_o = 32'h00000000 /* 0x7684 */;
                7586: data_o = 32'h00000000 /* 0x7688 */;
                7587: data_o = 32'h00000000 /* 0x768c */;
                7588: data_o = 32'h00000000 /* 0x7690 */;
                7589: data_o = 32'h00000000 /* 0x7694 */;
                7590: data_o = 32'h00000000 /* 0x7698 */;
                7591: data_o = 32'h00000000 /* 0x769c */;
                7592: data_o = 32'h00000000 /* 0x76a0 */;
                7593: data_o = 32'h00000000 /* 0x76a4 */;
                7594: data_o = 32'h00000000 /* 0x76a8 */;
                7595: data_o = 32'h00000000 /* 0x76ac */;
                7596: data_o = 32'h00000000 /* 0x76b0 */;
                7597: data_o = 32'h00000000 /* 0x76b4 */;
                7598: data_o = 32'h00000000 /* 0x76b8 */;
                7599: data_o = 32'h00000000 /* 0x76bc */;
                7600: data_o = 32'h00000000 /* 0x76c0 */;
                7601: data_o = 32'h00000000 /* 0x76c4 */;
                7602: data_o = 32'h00000000 /* 0x76c8 */;
                7603: data_o = 32'h00000000 /* 0x76cc */;
                7604: data_o = 32'h00000000 /* 0x76d0 */;
                7605: data_o = 32'h00000000 /* 0x76d4 */;
                7606: data_o = 32'h00000000 /* 0x76d8 */;
                7607: data_o = 32'h00000000 /* 0x76dc */;
                7608: data_o = 32'h00000000 /* 0x76e0 */;
                7609: data_o = 32'h00000000 /* 0x76e4 */;
                7610: data_o = 32'h00000000 /* 0x76e8 */;
                7611: data_o = 32'h00000000 /* 0x76ec */;
                7612: data_o = 32'h00000000 /* 0x76f0 */;
                7613: data_o = 32'h00000000 /* 0x76f4 */;
                7614: data_o = 32'h00000000 /* 0x76f8 */;
                7615: data_o = 32'h00000000 /* 0x76fc */;
                7616: data_o = 32'h00000000 /* 0x7700 */;
                7617: data_o = 32'h00000000 /* 0x7704 */;
                7618: data_o = 32'h00000000 /* 0x7708 */;
                7619: data_o = 32'h00000000 /* 0x770c */;
                7620: data_o = 32'h00000000 /* 0x7710 */;
                7621: data_o = 32'h00000000 /* 0x7714 */;
                7622: data_o = 32'h00000000 /* 0x7718 */;
                7623: data_o = 32'h00000000 /* 0x771c */;
                7624: data_o = 32'h00000000 /* 0x7720 */;
                7625: data_o = 32'h00000000 /* 0x7724 */;
                7626: data_o = 32'h00000000 /* 0x7728 */;
                7627: data_o = 32'h00000000 /* 0x772c */;
                7628: data_o = 32'h00000000 /* 0x7730 */;
                7629: data_o = 32'h00000000 /* 0x7734 */;
                7630: data_o = 32'h00000000 /* 0x7738 */;
                7631: data_o = 32'h00000000 /* 0x773c */;
                7632: data_o = 32'h00000000 /* 0x7740 */;
                7633: data_o = 32'h00000000 /* 0x7744 */;
                7634: data_o = 32'h00000000 /* 0x7748 */;
                7635: data_o = 32'h00000000 /* 0x774c */;
                7636: data_o = 32'h00000000 /* 0x7750 */;
                7637: data_o = 32'h00000000 /* 0x7754 */;
                7638: data_o = 32'h00000000 /* 0x7758 */;
                7639: data_o = 32'h00000000 /* 0x775c */;
                7640: data_o = 32'h00000000 /* 0x7760 */;
                7641: data_o = 32'h00000000 /* 0x7764 */;
                7642: data_o = 32'h00000000 /* 0x7768 */;
                7643: data_o = 32'h00000000 /* 0x776c */;
                7644: data_o = 32'h00000000 /* 0x7770 */;
                7645: data_o = 32'h00000000 /* 0x7774 */;
                7646: data_o = 32'h00000000 /* 0x7778 */;
                7647: data_o = 32'h00000000 /* 0x777c */;
                7648: data_o = 32'h00000000 /* 0x7780 */;
                7649: data_o = 32'h00000000 /* 0x7784 */;
                7650: data_o = 32'h00000000 /* 0x7788 */;
                7651: data_o = 32'h00000000 /* 0x778c */;
                7652: data_o = 32'h00000000 /* 0x7790 */;
                7653: data_o = 32'h00000000 /* 0x7794 */;
                7654: data_o = 32'h00000000 /* 0x7798 */;
                7655: data_o = 32'h00000000 /* 0x779c */;
                7656: data_o = 32'h00000000 /* 0x77a0 */;
                7657: data_o = 32'h00000000 /* 0x77a4 */;
                7658: data_o = 32'h00000000 /* 0x77a8 */;
                7659: data_o = 32'h00000000 /* 0x77ac */;
                7660: data_o = 32'h00000000 /* 0x77b0 */;
                7661: data_o = 32'h00000000 /* 0x77b4 */;
                7662: data_o = 32'h00000000 /* 0x77b8 */;
                7663: data_o = 32'h00000000 /* 0x77bc */;
                7664: data_o = 32'h00000000 /* 0x77c0 */;
                7665: data_o = 32'h00000000 /* 0x77c4 */;
                7666: data_o = 32'h00000000 /* 0x77c8 */;
                7667: data_o = 32'h00000000 /* 0x77cc */;
                7668: data_o = 32'h00000000 /* 0x77d0 */;
                7669: data_o = 32'h00000000 /* 0x77d4 */;
                7670: data_o = 32'h00000000 /* 0x77d8 */;
                7671: data_o = 32'h00000000 /* 0x77dc */;
                7672: data_o = 32'h00000000 /* 0x77e0 */;
                7673: data_o = 32'h00000000 /* 0x77e4 */;
                7674: data_o = 32'h00000000 /* 0x77e8 */;
                7675: data_o = 32'h00000000 /* 0x77ec */;
                7676: data_o = 32'h00000000 /* 0x77f0 */;
                7677: data_o = 32'h00000000 /* 0x77f4 */;
                7678: data_o = 32'h00000000 /* 0x77f8 */;
                7679: data_o = 32'h00000000 /* 0x77fc */;
                7680: data_o = 32'h00000000 /* 0x7800 */;
                7681: data_o = 32'h00000000 /* 0x7804 */;
                7682: data_o = 32'h00000000 /* 0x7808 */;
                7683: data_o = 32'h00000000 /* 0x780c */;
                7684: data_o = 32'h00000000 /* 0x7810 */;
                7685: data_o = 32'h00000000 /* 0x7814 */;
                7686: data_o = 32'h00000000 /* 0x7818 */;
                7687: data_o = 32'h00000000 /* 0x781c */;
                7688: data_o = 32'h00000000 /* 0x7820 */;
                7689: data_o = 32'h00000000 /* 0x7824 */;
                7690: data_o = 32'h00000000 /* 0x7828 */;
                7691: data_o = 32'h00000000 /* 0x782c */;
                7692: data_o = 32'h00000000 /* 0x7830 */;
                7693: data_o = 32'h00000000 /* 0x7834 */;
                7694: data_o = 32'h00000000 /* 0x7838 */;
                7695: data_o = 32'h00000000 /* 0x783c */;
                7696: data_o = 32'h00000000 /* 0x7840 */;
                7697: data_o = 32'h00000000 /* 0x7844 */;
                7698: data_o = 32'h00000000 /* 0x7848 */;
                7699: data_o = 32'h00000000 /* 0x784c */;
                7700: data_o = 32'h00000000 /* 0x7850 */;
                7701: data_o = 32'h00000000 /* 0x7854 */;
                7702: data_o = 32'h00000000 /* 0x7858 */;
                7703: data_o = 32'h00000000 /* 0x785c */;
                7704: data_o = 32'h00000000 /* 0x7860 */;
                7705: data_o = 32'h00000000 /* 0x7864 */;
                7706: data_o = 32'h00000000 /* 0x7868 */;
                7707: data_o = 32'h00000000 /* 0x786c */;
                7708: data_o = 32'h00000000 /* 0x7870 */;
                7709: data_o = 32'h00000000 /* 0x7874 */;
                7710: data_o = 32'h00000000 /* 0x7878 */;
                7711: data_o = 32'h00000000 /* 0x787c */;
                7712: data_o = 32'h00000000 /* 0x7880 */;
                7713: data_o = 32'h00000000 /* 0x7884 */;
                7714: data_o = 32'h00000000 /* 0x7888 */;
                7715: data_o = 32'h00000000 /* 0x788c */;
                7716: data_o = 32'h00000000 /* 0x7890 */;
                7717: data_o = 32'h00000000 /* 0x7894 */;
                7718: data_o = 32'h00000000 /* 0x7898 */;
                7719: data_o = 32'h00000000 /* 0x789c */;
                7720: data_o = 32'h00000000 /* 0x78a0 */;
                7721: data_o = 32'h00000000 /* 0x78a4 */;
                7722: data_o = 32'h00000000 /* 0x78a8 */;
                7723: data_o = 32'h00000000 /* 0x78ac */;
                7724: data_o = 32'h00000000 /* 0x78b0 */;
                7725: data_o = 32'h00000000 /* 0x78b4 */;
                7726: data_o = 32'h00000000 /* 0x78b8 */;
                7727: data_o = 32'h00000000 /* 0x78bc */;
                7728: data_o = 32'h00000000 /* 0x78c0 */;
                7729: data_o = 32'h00000000 /* 0x78c4 */;
                7730: data_o = 32'h00000000 /* 0x78c8 */;
                7731: data_o = 32'h00000000 /* 0x78cc */;
                7732: data_o = 32'h00000000 /* 0x78d0 */;
                7733: data_o = 32'h00000000 /* 0x78d4 */;
                7734: data_o = 32'h00000000 /* 0x78d8 */;
                7735: data_o = 32'h00000000 /* 0x78dc */;
                7736: data_o = 32'h00000000 /* 0x78e0 */;
                7737: data_o = 32'h00000000 /* 0x78e4 */;
                7738: data_o = 32'h00000000 /* 0x78e8 */;
                7739: data_o = 32'h00000000 /* 0x78ec */;
                7740: data_o = 32'h00000000 /* 0x78f0 */;
                7741: data_o = 32'h00000000 /* 0x78f4 */;
                7742: data_o = 32'h00000000 /* 0x78f8 */;
                7743: data_o = 32'h00000000 /* 0x78fc */;
                7744: data_o = 32'h00000000 /* 0x7900 */;
                7745: data_o = 32'h00000000 /* 0x7904 */;
                7746: data_o = 32'h00000000 /* 0x7908 */;
                7747: data_o = 32'h00000000 /* 0x790c */;
                7748: data_o = 32'h00000000 /* 0x7910 */;
                7749: data_o = 32'h00000000 /* 0x7914 */;
                7750: data_o = 32'h00000000 /* 0x7918 */;
                7751: data_o = 32'h00000000 /* 0x791c */;
                7752: data_o = 32'h00000000 /* 0x7920 */;
                7753: data_o = 32'h00000000 /* 0x7924 */;
                7754: data_o = 32'h00000000 /* 0x7928 */;
                7755: data_o = 32'h00000000 /* 0x792c */;
                7756: data_o = 32'h00000000 /* 0x7930 */;
                7757: data_o = 32'h00000000 /* 0x7934 */;
                7758: data_o = 32'h00000000 /* 0x7938 */;
                7759: data_o = 32'h00000000 /* 0x793c */;
                7760: data_o = 32'h00000000 /* 0x7940 */;
                7761: data_o = 32'h00000000 /* 0x7944 */;
                7762: data_o = 32'h00000000 /* 0x7948 */;
                7763: data_o = 32'h00000000 /* 0x794c */;
                7764: data_o = 32'h00000000 /* 0x7950 */;
                7765: data_o = 32'h00000000 /* 0x7954 */;
                7766: data_o = 32'h00000000 /* 0x7958 */;
                7767: data_o = 32'h00000000 /* 0x795c */;
                7768: data_o = 32'h00000000 /* 0x7960 */;
                7769: data_o = 32'h00000000 /* 0x7964 */;
                7770: data_o = 32'h00000000 /* 0x7968 */;
                7771: data_o = 32'h00000000 /* 0x796c */;
                7772: data_o = 32'h00000000 /* 0x7970 */;
                7773: data_o = 32'h00000000 /* 0x7974 */;
                7774: data_o = 32'h00000000 /* 0x7978 */;
                7775: data_o = 32'h00000000 /* 0x797c */;
                7776: data_o = 32'h00000000 /* 0x7980 */;
                7777: data_o = 32'h00000000 /* 0x7984 */;
                7778: data_o = 32'h00000000 /* 0x7988 */;
                7779: data_o = 32'h00000000 /* 0x798c */;
                7780: data_o = 32'h00000000 /* 0x7990 */;
                7781: data_o = 32'h00000000 /* 0x7994 */;
                7782: data_o = 32'h00000000 /* 0x7998 */;
                7783: data_o = 32'h00000000 /* 0x799c */;
                7784: data_o = 32'h00000000 /* 0x79a0 */;
                7785: data_o = 32'h00000000 /* 0x79a4 */;
                7786: data_o = 32'h00000000 /* 0x79a8 */;
                7787: data_o = 32'h00000000 /* 0x79ac */;
                7788: data_o = 32'h00000000 /* 0x79b0 */;
                7789: data_o = 32'h00000000 /* 0x79b4 */;
                7790: data_o = 32'h00000000 /* 0x79b8 */;
                7791: data_o = 32'h00000000 /* 0x79bc */;
                7792: data_o = 32'h00000000 /* 0x79c0 */;
                7793: data_o = 32'h00000000 /* 0x79c4 */;
                7794: data_o = 32'h00000000 /* 0x79c8 */;
                7795: data_o = 32'h00000000 /* 0x79cc */;
                7796: data_o = 32'h00000000 /* 0x79d0 */;
                7797: data_o = 32'h00000000 /* 0x79d4 */;
                7798: data_o = 32'h00000000 /* 0x79d8 */;
                7799: data_o = 32'h00000000 /* 0x79dc */;
                7800: data_o = 32'h00000000 /* 0x79e0 */;
                7801: data_o = 32'h00000000 /* 0x79e4 */;
                7802: data_o = 32'h00000000 /* 0x79e8 */;
                7803: data_o = 32'h00000000 /* 0x79ec */;
                7804: data_o = 32'h00000000 /* 0x79f0 */;
                7805: data_o = 32'h00000000 /* 0x79f4 */;
                7806: data_o = 32'h00000000 /* 0x79f8 */;
                7807: data_o = 32'h00000000 /* 0x79fc */;
                7808: data_o = 32'h00000000 /* 0x7a00 */;
                7809: data_o = 32'h00000000 /* 0x7a04 */;
                7810: data_o = 32'h00000000 /* 0x7a08 */;
                7811: data_o = 32'h00000000 /* 0x7a0c */;
                7812: data_o = 32'h00000000 /* 0x7a10 */;
                7813: data_o = 32'h00000000 /* 0x7a14 */;
                7814: data_o = 32'h00000000 /* 0x7a18 */;
                7815: data_o = 32'h00000000 /* 0x7a1c */;
                7816: data_o = 32'h00000000 /* 0x7a20 */;
                7817: data_o = 32'h00000000 /* 0x7a24 */;
                7818: data_o = 32'h00000000 /* 0x7a28 */;
                7819: data_o = 32'h00000000 /* 0x7a2c */;
                7820: data_o = 32'h00000000 /* 0x7a30 */;
                7821: data_o = 32'h00000000 /* 0x7a34 */;
                7822: data_o = 32'h00000000 /* 0x7a38 */;
                7823: data_o = 32'h00000000 /* 0x7a3c */;
                7824: data_o = 32'h00000000 /* 0x7a40 */;
                7825: data_o = 32'h00000000 /* 0x7a44 */;
                7826: data_o = 32'h00000000 /* 0x7a48 */;
                7827: data_o = 32'h00000000 /* 0x7a4c */;
                7828: data_o = 32'h00000000 /* 0x7a50 */;
                7829: data_o = 32'h00000000 /* 0x7a54 */;
                7830: data_o = 32'h00000000 /* 0x7a58 */;
                7831: data_o = 32'h00000000 /* 0x7a5c */;
                7832: data_o = 32'h00000000 /* 0x7a60 */;
                7833: data_o = 32'h00000000 /* 0x7a64 */;
                7834: data_o = 32'h00000000 /* 0x7a68 */;
                7835: data_o = 32'h00000000 /* 0x7a6c */;
                7836: data_o = 32'h00000000 /* 0x7a70 */;
                7837: data_o = 32'h00000000 /* 0x7a74 */;
                7838: data_o = 32'h00000000 /* 0x7a78 */;
                7839: data_o = 32'h00000000 /* 0x7a7c */;
                7840: data_o = 32'h00000000 /* 0x7a80 */;
                7841: data_o = 32'h00000000 /* 0x7a84 */;
                7842: data_o = 32'h00000000 /* 0x7a88 */;
                7843: data_o = 32'h00000000 /* 0x7a8c */;
                7844: data_o = 32'h00000000 /* 0x7a90 */;
                7845: data_o = 32'h00000000 /* 0x7a94 */;
                7846: data_o = 32'h00000000 /* 0x7a98 */;
                7847: data_o = 32'h00000000 /* 0x7a9c */;
                7848: data_o = 32'h00000000 /* 0x7aa0 */;
                7849: data_o = 32'h00000000 /* 0x7aa4 */;
                7850: data_o = 32'h00000000 /* 0x7aa8 */;
                7851: data_o = 32'h00000000 /* 0x7aac */;
                7852: data_o = 32'h00000000 /* 0x7ab0 */;
                7853: data_o = 32'h00000000 /* 0x7ab4 */;
                7854: data_o = 32'h00000000 /* 0x7ab8 */;
                7855: data_o = 32'h00000000 /* 0x7abc */;
                7856: data_o = 32'h00000000 /* 0x7ac0 */;
                7857: data_o = 32'h00000000 /* 0x7ac4 */;
                7858: data_o = 32'h00000000 /* 0x7ac8 */;
                7859: data_o = 32'h00000000 /* 0x7acc */;
                7860: data_o = 32'h00000000 /* 0x7ad0 */;
                7861: data_o = 32'h00000000 /* 0x7ad4 */;
                7862: data_o = 32'h00000000 /* 0x7ad8 */;
                7863: data_o = 32'h00000000 /* 0x7adc */;
                7864: data_o = 32'h00000000 /* 0x7ae0 */;
                7865: data_o = 32'h00000000 /* 0x7ae4 */;
                7866: data_o = 32'h00000000 /* 0x7ae8 */;
                7867: data_o = 32'h00000000 /* 0x7aec */;
                7868: data_o = 32'h00000000 /* 0x7af0 */;
                7869: data_o = 32'h00000000 /* 0x7af4 */;
                7870: data_o = 32'h00000000 /* 0x7af8 */;
                7871: data_o = 32'h00000000 /* 0x7afc */;
                7872: data_o = 32'h00000000 /* 0x7b00 */;
                7873: data_o = 32'h00000000 /* 0x7b04 */;
                7874: data_o = 32'h00000000 /* 0x7b08 */;
                7875: data_o = 32'h00000000 /* 0x7b0c */;
                7876: data_o = 32'h00000000 /* 0x7b10 */;
                7877: data_o = 32'h00000000 /* 0x7b14 */;
                7878: data_o = 32'h00000000 /* 0x7b18 */;
                7879: data_o = 32'h00000000 /* 0x7b1c */;
                7880: data_o = 32'h00000000 /* 0x7b20 */;
                7881: data_o = 32'h00000000 /* 0x7b24 */;
                7882: data_o = 32'h00000000 /* 0x7b28 */;
                7883: data_o = 32'h00000000 /* 0x7b2c */;
                7884: data_o = 32'h00000000 /* 0x7b30 */;
                7885: data_o = 32'h00000000 /* 0x7b34 */;
                7886: data_o = 32'h00000000 /* 0x7b38 */;
                7887: data_o = 32'h00000000 /* 0x7b3c */;
                7888: data_o = 32'h00000000 /* 0x7b40 */;
                7889: data_o = 32'h00000000 /* 0x7b44 */;
                7890: data_o = 32'h00000000 /* 0x7b48 */;
                7891: data_o = 32'h00000000 /* 0x7b4c */;
                7892: data_o = 32'h00000000 /* 0x7b50 */;
                7893: data_o = 32'h00000000 /* 0x7b54 */;
                7894: data_o = 32'h00000000 /* 0x7b58 */;
                7895: data_o = 32'h00000000 /* 0x7b5c */;
                7896: data_o = 32'h00000000 /* 0x7b60 */;
                7897: data_o = 32'h00000000 /* 0x7b64 */;
                7898: data_o = 32'h00000000 /* 0x7b68 */;
                7899: data_o = 32'h00000000 /* 0x7b6c */;
                7900: data_o = 32'h00000000 /* 0x7b70 */;
                7901: data_o = 32'h00000000 /* 0x7b74 */;
                7902: data_o = 32'h00000000 /* 0x7b78 */;
                7903: data_o = 32'h00000000 /* 0x7b7c */;
                7904: data_o = 32'h00000000 /* 0x7b80 */;
                7905: data_o = 32'h00000000 /* 0x7b84 */;
                7906: data_o = 32'h00000000 /* 0x7b88 */;
                7907: data_o = 32'h00000000 /* 0x7b8c */;
                7908: data_o = 32'h00000000 /* 0x7b90 */;
                7909: data_o = 32'h00000000 /* 0x7b94 */;
                7910: data_o = 32'h00000000 /* 0x7b98 */;
                7911: data_o = 32'h00000000 /* 0x7b9c */;
                7912: data_o = 32'h00000000 /* 0x7ba0 */;
                7913: data_o = 32'h00000000 /* 0x7ba4 */;
                7914: data_o = 32'h00000000 /* 0x7ba8 */;
                7915: data_o = 32'h00000000 /* 0x7bac */;
                7916: data_o = 32'h00000000 /* 0x7bb0 */;
                7917: data_o = 32'h00000000 /* 0x7bb4 */;
                7918: data_o = 32'h00000000 /* 0x7bb8 */;
                7919: data_o = 32'h00000000 /* 0x7bbc */;
                7920: data_o = 32'h00000000 /* 0x7bc0 */;
                7921: data_o = 32'h00000000 /* 0x7bc4 */;
                7922: data_o = 32'h00000000 /* 0x7bc8 */;
                7923: data_o = 32'h00000000 /* 0x7bcc */;
                7924: data_o = 32'h00000000 /* 0x7bd0 */;
                7925: data_o = 32'h00000000 /* 0x7bd4 */;
                7926: data_o = 32'h00000000 /* 0x7bd8 */;
                7927: data_o = 32'h00000000 /* 0x7bdc */;
                7928: data_o = 32'h00000000 /* 0x7be0 */;
                7929: data_o = 32'h00000000 /* 0x7be4 */;
                7930: data_o = 32'h00000000 /* 0x7be8 */;
                7931: data_o = 32'h00000000 /* 0x7bec */;
                7932: data_o = 32'h00000000 /* 0x7bf0 */;
                7933: data_o = 32'h00000000 /* 0x7bf4 */;
                7934: data_o = 32'h00000000 /* 0x7bf8 */;
                7935: data_o = 32'h00000000 /* 0x7bfc */;
                7936: data_o = 32'h00000000 /* 0x7c00 */;
                7937: data_o = 32'h00000000 /* 0x7c04 */;
                7938: data_o = 32'h00000000 /* 0x7c08 */;
                7939: data_o = 32'h00000000 /* 0x7c0c */;
                7940: data_o = 32'h00000000 /* 0x7c10 */;
                7941: data_o = 32'h00000000 /* 0x7c14 */;
                7942: data_o = 32'h00000000 /* 0x7c18 */;
                7943: data_o = 32'h00000000 /* 0x7c1c */;
                7944: data_o = 32'h00000000 /* 0x7c20 */;
                7945: data_o = 32'h00000000 /* 0x7c24 */;
                7946: data_o = 32'h00000000 /* 0x7c28 */;
                7947: data_o = 32'h00000000 /* 0x7c2c */;
                7948: data_o = 32'h00000000 /* 0x7c30 */;
                7949: data_o = 32'h00000000 /* 0x7c34 */;
                7950: data_o = 32'h00000000 /* 0x7c38 */;
                7951: data_o = 32'h00000000 /* 0x7c3c */;
                7952: data_o = 32'h00000000 /* 0x7c40 */;
                7953: data_o = 32'h00000000 /* 0x7c44 */;
                7954: data_o = 32'h00000000 /* 0x7c48 */;
                7955: data_o = 32'h00000000 /* 0x7c4c */;
                7956: data_o = 32'h00000000 /* 0x7c50 */;
                7957: data_o = 32'h00000000 /* 0x7c54 */;
                7958: data_o = 32'h00000000 /* 0x7c58 */;
                7959: data_o = 32'h00000000 /* 0x7c5c */;
                7960: data_o = 32'h00000000 /* 0x7c60 */;
                7961: data_o = 32'h00000000 /* 0x7c64 */;
                7962: data_o = 32'h00000000 /* 0x7c68 */;
                7963: data_o = 32'h00000000 /* 0x7c6c */;
                7964: data_o = 32'h00000000 /* 0x7c70 */;
                7965: data_o = 32'h00000000 /* 0x7c74 */;
                7966: data_o = 32'h00000000 /* 0x7c78 */;
                7967: data_o = 32'h00000000 /* 0x7c7c */;
                7968: data_o = 32'h00000000 /* 0x7c80 */;
                7969: data_o = 32'h00000000 /* 0x7c84 */;
                7970: data_o = 32'h00000000 /* 0x7c88 */;
                7971: data_o = 32'h00000000 /* 0x7c8c */;
                7972: data_o = 32'h00000000 /* 0x7c90 */;
                7973: data_o = 32'h00000000 /* 0x7c94 */;
                7974: data_o = 32'h00000000 /* 0x7c98 */;
                7975: data_o = 32'h00000000 /* 0x7c9c */;
                7976: data_o = 32'h00000000 /* 0x7ca0 */;
                7977: data_o = 32'h00000000 /* 0x7ca4 */;
                7978: data_o = 32'h00000000 /* 0x7ca8 */;
                7979: data_o = 32'h00000000 /* 0x7cac */;
                7980: data_o = 32'h00000000 /* 0x7cb0 */;
                7981: data_o = 32'h00000000 /* 0x7cb4 */;
                7982: data_o = 32'h00000000 /* 0x7cb8 */;
                7983: data_o = 32'h00000000 /* 0x7cbc */;
                7984: data_o = 32'h00000000 /* 0x7cc0 */;
                7985: data_o = 32'h00000000 /* 0x7cc4 */;
                7986: data_o = 32'h00000000 /* 0x7cc8 */;
                7987: data_o = 32'h00000000 /* 0x7ccc */;
                7988: data_o = 32'h00000000 /* 0x7cd0 */;
                7989: data_o = 32'h00000000 /* 0x7cd4 */;
                7990: data_o = 32'h00000000 /* 0x7cd8 */;
                7991: data_o = 32'h00000000 /* 0x7cdc */;
                7992: data_o = 32'h00000000 /* 0x7ce0 */;
                7993: data_o = 32'h00000000 /* 0x7ce4 */;
                7994: data_o = 32'h00000000 /* 0x7ce8 */;
                7995: data_o = 32'h00000000 /* 0x7cec */;
                7996: data_o = 32'h00000000 /* 0x7cf0 */;
                7997: data_o = 32'h00000000 /* 0x7cf4 */;
                7998: data_o = 32'h00000000 /* 0x7cf8 */;
                7999: data_o = 32'h00000000 /* 0x7cfc */;
                8000: data_o = 32'h00000000 /* 0x7d00 */;
                8001: data_o = 32'h00000000 /* 0x7d04 */;
                8002: data_o = 32'h00000000 /* 0x7d08 */;
                8003: data_o = 32'h00000000 /* 0x7d0c */;
                8004: data_o = 32'h00000000 /* 0x7d10 */;
                8005: data_o = 32'h00000000 /* 0x7d14 */;
                8006: data_o = 32'h00000000 /* 0x7d18 */;
                8007: data_o = 32'h00000000 /* 0x7d1c */;
                8008: data_o = 32'h00000000 /* 0x7d20 */;
                8009: data_o = 32'h00000000 /* 0x7d24 */;
                8010: data_o = 32'h00000000 /* 0x7d28 */;
                8011: data_o = 32'h00000000 /* 0x7d2c */;
                8012: data_o = 32'h00000000 /* 0x7d30 */;
                8013: data_o = 32'h00000000 /* 0x7d34 */;
                8014: data_o = 32'h00000000 /* 0x7d38 */;
                8015: data_o = 32'h00000000 /* 0x7d3c */;
                8016: data_o = 32'h00000000 /* 0x7d40 */;
                8017: data_o = 32'h00000000 /* 0x7d44 */;
                8018: data_o = 32'h00000000 /* 0x7d48 */;
                8019: data_o = 32'h00000000 /* 0x7d4c */;
                8020: data_o = 32'h00000000 /* 0x7d50 */;
                8021: data_o = 32'h00000000 /* 0x7d54 */;
                8022: data_o = 32'h00000000 /* 0x7d58 */;
                8023: data_o = 32'h00000000 /* 0x7d5c */;
                8024: data_o = 32'h00000000 /* 0x7d60 */;
                8025: data_o = 32'h00000000 /* 0x7d64 */;
                8026: data_o = 32'h00000000 /* 0x7d68 */;
                8027: data_o = 32'h00000000 /* 0x7d6c */;
                8028: data_o = 32'h00000000 /* 0x7d70 */;
                8029: data_o = 32'h00000000 /* 0x7d74 */;
                8030: data_o = 32'h00000000 /* 0x7d78 */;
                8031: data_o = 32'h00000000 /* 0x7d7c */;
                8032: data_o = 32'h00000000 /* 0x7d80 */;
                8033: data_o = 32'h00000000 /* 0x7d84 */;
                8034: data_o = 32'h00000000 /* 0x7d88 */;
                8035: data_o = 32'h00000000 /* 0x7d8c */;
                8036: data_o = 32'h00000000 /* 0x7d90 */;
                8037: data_o = 32'h00000000 /* 0x7d94 */;
                8038: data_o = 32'h00000000 /* 0x7d98 */;
                8039: data_o = 32'h00000000 /* 0x7d9c */;
                8040: data_o = 32'h00000000 /* 0x7da0 */;
                8041: data_o = 32'h00000000 /* 0x7da4 */;
                8042: data_o = 32'h00000000 /* 0x7da8 */;
                8043: data_o = 32'h00000000 /* 0x7dac */;
                8044: data_o = 32'h00000000 /* 0x7db0 */;
                8045: data_o = 32'h00000000 /* 0x7db4 */;
                8046: data_o = 32'h00000000 /* 0x7db8 */;
                8047: data_o = 32'h00000000 /* 0x7dbc */;
                8048: data_o = 32'h00000000 /* 0x7dc0 */;
                8049: data_o = 32'h00000000 /* 0x7dc4 */;
                8050: data_o = 32'h00000000 /* 0x7dc8 */;
                8051: data_o = 32'h00000000 /* 0x7dcc */;
                8052: data_o = 32'h00000000 /* 0x7dd0 */;
                8053: data_o = 32'h00000000 /* 0x7dd4 */;
                8054: data_o = 32'h00000000 /* 0x7dd8 */;
                8055: data_o = 32'h00000000 /* 0x7ddc */;
                8056: data_o = 32'h00000000 /* 0x7de0 */;
                8057: data_o = 32'h00000000 /* 0x7de4 */;
                8058: data_o = 32'h00000000 /* 0x7de8 */;
                8059: data_o = 32'h00000000 /* 0x7dec */;
                8060: data_o = 32'h00000000 /* 0x7df0 */;
                8061: data_o = 32'h00000000 /* 0x7df4 */;
                8062: data_o = 32'h00000000 /* 0x7df8 */;
                8063: data_o = 32'h00000000 /* 0x7dfc */;
                8064: data_o = 32'h00000000 /* 0x7e00 */;
                8065: data_o = 32'h00000000 /* 0x7e04 */;
                8066: data_o = 32'h00000000 /* 0x7e08 */;
                8067: data_o = 32'h00000000 /* 0x7e0c */;
                8068: data_o = 32'h00000000 /* 0x7e10 */;
                8069: data_o = 32'h00000000 /* 0x7e14 */;
                8070: data_o = 32'h00000000 /* 0x7e18 */;
                8071: data_o = 32'h00000000 /* 0x7e1c */;
                8072: data_o = 32'h00000000 /* 0x7e20 */;
                8073: data_o = 32'h00000000 /* 0x7e24 */;
                8074: data_o = 32'h00000000 /* 0x7e28 */;
                8075: data_o = 32'h00000000 /* 0x7e2c */;
                8076: data_o = 32'h00000000 /* 0x7e30 */;
                8077: data_o = 32'h00000000 /* 0x7e34 */;
                8078: data_o = 32'h00000000 /* 0x7e38 */;
                8079: data_o = 32'h00000000 /* 0x7e3c */;
                8080: data_o = 32'h00000000 /* 0x7e40 */;
                8081: data_o = 32'h00000000 /* 0x7e44 */;
                8082: data_o = 32'h00000000 /* 0x7e48 */;
                8083: data_o = 32'h00000000 /* 0x7e4c */;
                8084: data_o = 32'h00000000 /* 0x7e50 */;
                8085: data_o = 32'h00000000 /* 0x7e54 */;
                8086: data_o = 32'h00000000 /* 0x7e58 */;
                8087: data_o = 32'h00000000 /* 0x7e5c */;
                8088: data_o = 32'h00000000 /* 0x7e60 */;
                8089: data_o = 32'h00000000 /* 0x7e64 */;
                8090: data_o = 32'h00000000 /* 0x7e68 */;
                8091: data_o = 32'h00000000 /* 0x7e6c */;
                8092: data_o = 32'h00000000 /* 0x7e70 */;
                8093: data_o = 32'h00000000 /* 0x7e74 */;
                8094: data_o = 32'h00000000 /* 0x7e78 */;
                8095: data_o = 32'h00000000 /* 0x7e7c */;
                8096: data_o = 32'h00000000 /* 0x7e80 */;
                8097: data_o = 32'h00000000 /* 0x7e84 */;
                8098: data_o = 32'h00000000 /* 0x7e88 */;
                8099: data_o = 32'h00000000 /* 0x7e8c */;
                8100: data_o = 32'h00000000 /* 0x7e90 */;
                8101: data_o = 32'h00000000 /* 0x7e94 */;
                8102: data_o = 32'h00000000 /* 0x7e98 */;
                8103: data_o = 32'h00000000 /* 0x7e9c */;
                8104: data_o = 32'h00000000 /* 0x7ea0 */;
                8105: data_o = 32'h00000000 /* 0x7ea4 */;
                8106: data_o = 32'h00000000 /* 0x7ea8 */;
                8107: data_o = 32'h00000000 /* 0x7eac */;
                8108: data_o = 32'h00000000 /* 0x7eb0 */;
                8109: data_o = 32'h00000000 /* 0x7eb4 */;
                8110: data_o = 32'h00000000 /* 0x7eb8 */;
                8111: data_o = 32'h00000000 /* 0x7ebc */;
                8112: data_o = 32'h00000000 /* 0x7ec0 */;
                8113: data_o = 32'h00000000 /* 0x7ec4 */;
                8114: data_o = 32'h00000000 /* 0x7ec8 */;
                8115: data_o = 32'h00000000 /* 0x7ecc */;
                8116: data_o = 32'h00000000 /* 0x7ed0 */;
                8117: data_o = 32'h00000000 /* 0x7ed4 */;
                8118: data_o = 32'h00000000 /* 0x7ed8 */;
                8119: data_o = 32'h00000000 /* 0x7edc */;
                8120: data_o = 32'h00000000 /* 0x7ee0 */;
                8121: data_o = 32'h00000000 /* 0x7ee4 */;
                8122: data_o = 32'h00000000 /* 0x7ee8 */;
                8123: data_o = 32'h00000000 /* 0x7eec */;
                8124: data_o = 32'h00000000 /* 0x7ef0 */;
                8125: data_o = 32'h00000000 /* 0x7ef4 */;
                8126: data_o = 32'h00000000 /* 0x7ef8 */;
                8127: data_o = 32'h00000000 /* 0x7efc */;
                8128: data_o = 32'h00000000 /* 0x7f00 */;
                8129: data_o = 32'h00000000 /* 0x7f04 */;
                8130: data_o = 32'h00000000 /* 0x7f08 */;
                8131: data_o = 32'h00000000 /* 0x7f0c */;
                8132: data_o = 32'h00000000 /* 0x7f10 */;
                8133: data_o = 32'h00000000 /* 0x7f14 */;
                8134: data_o = 32'h00000000 /* 0x7f18 */;
                8135: data_o = 32'h00000000 /* 0x7f1c */;
                8136: data_o = 32'h00000000 /* 0x7f20 */;
                8137: data_o = 32'h00000000 /* 0x7f24 */;
                8138: data_o = 32'h00000000 /* 0x7f28 */;
                8139: data_o = 32'h00000000 /* 0x7f2c */;
                8140: data_o = 32'h00000000 /* 0x7f30 */;
                8141: data_o = 32'h00000000 /* 0x7f34 */;
                8142: data_o = 32'h00000000 /* 0x7f38 */;
                8143: data_o = 32'h00000000 /* 0x7f3c */;
                8144: data_o = 32'h00000000 /* 0x7f40 */;
                8145: data_o = 32'h00000000 /* 0x7f44 */;
                8146: data_o = 32'h00000000 /* 0x7f48 */;
                8147: data_o = 32'h00000000 /* 0x7f4c */;
                8148: data_o = 32'h00000000 /* 0x7f50 */;
                8149: data_o = 32'h00000000 /* 0x7f54 */;
                8150: data_o = 32'h00000000 /* 0x7f58 */;
                8151: data_o = 32'h00000000 /* 0x7f5c */;
                8152: data_o = 32'h00000000 /* 0x7f60 */;
                8153: data_o = 32'h00000000 /* 0x7f64 */;
                8154: data_o = 32'h00000000 /* 0x7f68 */;
                8155: data_o = 32'h00000000 /* 0x7f6c */;
                8156: data_o = 32'h00000000 /* 0x7f70 */;
                8157: data_o = 32'h00000000 /* 0x7f74 */;
                8158: data_o = 32'h00000000 /* 0x7f78 */;
                8159: data_o = 32'h00000000 /* 0x7f7c */;
                8160: data_o = 32'h00000000 /* 0x7f80 */;
                8161: data_o = 32'h00000000 /* 0x7f84 */;
                8162: data_o = 32'h00000000 /* 0x7f88 */;
                8163: data_o = 32'h00000000 /* 0x7f8c */;
                8164: data_o = 32'h00000000 /* 0x7f90 */;
                8165: data_o = 32'h00000000 /* 0x7f94 */;
                8166: data_o = 32'h00000000 /* 0x7f98 */;
                8167: data_o = 32'h00000000 /* 0x7f9c */;
                8168: data_o = 32'h00000000 /* 0x7fa0 */;
                8169: data_o = 32'h00000000 /* 0x7fa4 */;
                8170: data_o = 32'h00000000 /* 0x7fa8 */;
                8171: data_o = 32'h00000000 /* 0x7fac */;
                8172: data_o = 32'h00000000 /* 0x7fb0 */;
                8173: data_o = 32'h00000000 /* 0x7fb4 */;
                8174: data_o = 32'h00000000 /* 0x7fb8 */;
                8175: data_o = 32'h00000000 /* 0x7fbc */;
                8176: data_o = 32'h00000000 /* 0x7fc0 */;
                8177: data_o = 32'h00000000 /* 0x7fc4 */;
                8178: data_o = 32'h00000000 /* 0x7fc8 */;
                8179: data_o = 32'h00000000 /* 0x7fcc */;
                8180: data_o = 32'h00000000 /* 0x7fd0 */;
                8181: data_o = 32'h00000000 /* 0x7fd4 */;
                8182: data_o = 32'h00000000 /* 0x7fd8 */;
                8183: data_o = 32'h00000000 /* 0x7fdc */;
                8184: data_o = 32'h00000000 /* 0x7fe0 */;
                8185: data_o = 32'h00000000 /* 0x7fe4 */;
                8186: data_o = 32'h00000000 /* 0x7fe8 */;
                8187: data_o = 32'h00000000 /* 0x7fec */;
                8188: data_o = 32'h00000000 /* 0x7ff0 */;
                8189: data_o = 32'h00000000 /* 0x7ff4 */;
                8190: data_o = 32'h00000000 /* 0x7ff8 */;
                8191: data_o = 32'h00000000 /* 0x7ffc */;
                8192: data_o = 32'h00000000 /* 0x8000 */;
                8193: data_o = 32'h00000000 /* 0x8004 */;
                8194: data_o = 32'h00000000 /* 0x8008 */;
                8195: data_o = 32'h00000000 /* 0x800c */;
                8196: data_o = 32'h00000000 /* 0x8010 */;
                8197: data_o = 32'h00000000 /* 0x8014 */;
                8198: data_o = 32'h00000000 /* 0x8018 */;
                8199: data_o = 32'h00000000 /* 0x801c */;
                8200: data_o = 32'h00000000 /* 0x8020 */;
                8201: data_o = 32'h00000000 /* 0x8024 */;
                8202: data_o = 32'h00000000 /* 0x8028 */;
                8203: data_o = 32'h00000000 /* 0x802c */;
                8204: data_o = 32'h00000000 /* 0x8030 */;
                8205: data_o = 32'h00000000 /* 0x8034 */;
                8206: data_o = 32'h00000000 /* 0x8038 */;
                8207: data_o = 32'h00000000 /* 0x803c */;
                8208: data_o = 32'h00000000 /* 0x8040 */;
                8209: data_o = 32'h00000000 /* 0x8044 */;
                8210: data_o = 32'h00000000 /* 0x8048 */;
                8211: data_o = 32'h00000000 /* 0x804c */;
                8212: data_o = 32'h00000000 /* 0x8050 */;
                8213: data_o = 32'h00000000 /* 0x8054 */;
                8214: data_o = 32'h00000000 /* 0x8058 */;
                8215: data_o = 32'h00000000 /* 0x805c */;
                8216: data_o = 32'h00000000 /* 0x8060 */;
                8217: data_o = 32'h00000000 /* 0x8064 */;
                8218: data_o = 32'h00000000 /* 0x8068 */;
                8219: data_o = 32'h00000000 /* 0x806c */;
                8220: data_o = 32'h00000000 /* 0x8070 */;
                8221: data_o = 32'h00000000 /* 0x8074 */;
                8222: data_o = 32'h00000000 /* 0x8078 */;
                8223: data_o = 32'h00000000 /* 0x807c */;
                8224: data_o = 32'h00000000 /* 0x8080 */;
                8225: data_o = 32'h00000000 /* 0x8084 */;
                8226: data_o = 32'h00000000 /* 0x8088 */;
                8227: data_o = 32'h00000000 /* 0x808c */;
                8228: data_o = 32'h00000000 /* 0x8090 */;
                8229: data_o = 32'h00000000 /* 0x8094 */;
                8230: data_o = 32'h00000000 /* 0x8098 */;
                8231: data_o = 32'h00000000 /* 0x809c */;
                8232: data_o = 32'h00000000 /* 0x80a0 */;
                8233: data_o = 32'h00000000 /* 0x80a4 */;
                8234: data_o = 32'h00000000 /* 0x80a8 */;
                8235: data_o = 32'h00000000 /* 0x80ac */;
                8236: data_o = 32'h00000000 /* 0x80b0 */;
                8237: data_o = 32'h00000000 /* 0x80b4 */;
                8238: data_o = 32'h00000000 /* 0x80b8 */;
                8239: data_o = 32'h00000000 /* 0x80bc */;
                8240: data_o = 32'h00000000 /* 0x80c0 */;
                8241: data_o = 32'h00000000 /* 0x80c4 */;
                8242: data_o = 32'h00000000 /* 0x80c8 */;
                8243: data_o = 32'h00000000 /* 0x80cc */;
                8244: data_o = 32'h00000000 /* 0x80d0 */;
                8245: data_o = 32'h00000000 /* 0x80d4 */;
                8246: data_o = 32'h00000000 /* 0x80d8 */;
                8247: data_o = 32'h00000000 /* 0x80dc */;
                8248: data_o = 32'h00000000 /* 0x80e0 */;
                8249: data_o = 32'h00000000 /* 0x80e4 */;
                8250: data_o = 32'h00000000 /* 0x80e8 */;
                8251: data_o = 32'h00000000 /* 0x80ec */;
                8252: data_o = 32'h00000000 /* 0x80f0 */;
                8253: data_o = 32'h00000000 /* 0x80f4 */;
                8254: data_o = 32'h00000000 /* 0x80f8 */;
                8255: data_o = 32'h00000000 /* 0x80fc */;
                8256: data_o = 32'h00000000 /* 0x8100 */;
                8257: data_o = 32'h00000000 /* 0x8104 */;
                8258: data_o = 32'h00000000 /* 0x8108 */;
                8259: data_o = 32'h00000000 /* 0x810c */;
                8260: data_o = 32'h00000000 /* 0x8110 */;
                8261: data_o = 32'h00000000 /* 0x8114 */;
                8262: data_o = 32'h00000000 /* 0x8118 */;
                8263: data_o = 32'h00000000 /* 0x811c */;
                8264: data_o = 32'h00000000 /* 0x8120 */;
                8265: data_o = 32'h00000000 /* 0x8124 */;
                8266: data_o = 32'h00000000 /* 0x8128 */;
                8267: data_o = 32'h00000000 /* 0x812c */;
                8268: data_o = 32'h00000000 /* 0x8130 */;
                8269: data_o = 32'h00000000 /* 0x8134 */;
                8270: data_o = 32'h00000000 /* 0x8138 */;
                8271: data_o = 32'h00000000 /* 0x813c */;
                8272: data_o = 32'h00000000 /* 0x8140 */;
                8273: data_o = 32'h00000000 /* 0x8144 */;
                8274: data_o = 32'h00000000 /* 0x8148 */;
                8275: data_o = 32'h00000000 /* 0x814c */;
                8276: data_o = 32'h00000000 /* 0x8150 */;
                8277: data_o = 32'h00000000 /* 0x8154 */;
                8278: data_o = 32'h00000000 /* 0x8158 */;
                8279: data_o = 32'h00000000 /* 0x815c */;
                8280: data_o = 32'h00000000 /* 0x8160 */;
                8281: data_o = 32'h00000000 /* 0x8164 */;
                8282: data_o = 32'h00000000 /* 0x8168 */;
                8283: data_o = 32'h00000000 /* 0x816c */;
                8284: data_o = 32'h00000000 /* 0x8170 */;
                8285: data_o = 32'h00000000 /* 0x8174 */;
                8286: data_o = 32'h00000000 /* 0x8178 */;
                8287: data_o = 32'h00000000 /* 0x817c */;
                8288: data_o = 32'h00000000 /* 0x8180 */;
                8289: data_o = 32'h00000000 /* 0x8184 */;
                8290: data_o = 32'h00000000 /* 0x8188 */;
                8291: data_o = 32'h00000000 /* 0x818c */;
                8292: data_o = 32'h00000000 /* 0x8190 */;
                8293: data_o = 32'h00000000 /* 0x8194 */;
                8294: data_o = 32'h00000000 /* 0x8198 */;
                8295: data_o = 32'h00000000 /* 0x819c */;
                8296: data_o = 32'h00000000 /* 0x81a0 */;
                8297: data_o = 32'h00000000 /* 0x81a4 */;
                8298: data_o = 32'h00000000 /* 0x81a8 */;
                8299: data_o = 32'h00000000 /* 0x81ac */;
                8300: data_o = 32'h00000000 /* 0x81b0 */;
                8301: data_o = 32'h00000000 /* 0x81b4 */;
                8302: data_o = 32'h00000000 /* 0x81b8 */;
                8303: data_o = 32'h00000000 /* 0x81bc */;
                8304: data_o = 32'h00000000 /* 0x81c0 */;
                8305: data_o = 32'h00000000 /* 0x81c4 */;
                8306: data_o = 32'h00000000 /* 0x81c8 */;
                8307: data_o = 32'h00000000 /* 0x81cc */;
                8308: data_o = 32'h00000000 /* 0x81d0 */;
                8309: data_o = 32'h00000000 /* 0x81d4 */;
                8310: data_o = 32'h00000000 /* 0x81d8 */;
                8311: data_o = 32'h00000000 /* 0x81dc */;
                8312: data_o = 32'h00000000 /* 0x81e0 */;
                8313: data_o = 32'h00000000 /* 0x81e4 */;
                8314: data_o = 32'h00000000 /* 0x81e8 */;
                8315: data_o = 32'h00000000 /* 0x81ec */;
                8316: data_o = 32'h00000000 /* 0x81f0 */;
                8317: data_o = 32'h00000000 /* 0x81f4 */;
                8318: data_o = 32'h00000000 /* 0x81f8 */;
                8319: data_o = 32'h00000000 /* 0x81fc */;
                8320: data_o = 32'h00000000 /* 0x8200 */;
                8321: data_o = 32'h00000000 /* 0x8204 */;
                8322: data_o = 32'h00000000 /* 0x8208 */;
                8323: data_o = 32'h00000000 /* 0x820c */;
                8324: data_o = 32'h00000000 /* 0x8210 */;
                8325: data_o = 32'h00000000 /* 0x8214 */;
                8326: data_o = 32'h00000000 /* 0x8218 */;
                8327: data_o = 32'h00000000 /* 0x821c */;
                8328: data_o = 32'h00000000 /* 0x8220 */;
                8329: data_o = 32'h00000000 /* 0x8224 */;
                8330: data_o = 32'h00000000 /* 0x8228 */;
                8331: data_o = 32'h00000000 /* 0x822c */;
                8332: data_o = 32'h00000000 /* 0x8230 */;
                8333: data_o = 32'h00000000 /* 0x8234 */;
                8334: data_o = 32'h00000000 /* 0x8238 */;
                8335: data_o = 32'h00000000 /* 0x823c */;
                8336: data_o = 32'h00000000 /* 0x8240 */;
                8337: data_o = 32'h00000000 /* 0x8244 */;
                8338: data_o = 32'h00000000 /* 0x8248 */;
                8339: data_o = 32'h00000000 /* 0x824c */;
                8340: data_o = 32'h00000000 /* 0x8250 */;
                8341: data_o = 32'h00000000 /* 0x8254 */;
                8342: data_o = 32'h00000000 /* 0x8258 */;
                8343: data_o = 32'h00000000 /* 0x825c */;
                8344: data_o = 32'h00000000 /* 0x8260 */;
                8345: data_o = 32'h00000000 /* 0x8264 */;
                8346: data_o = 32'h00000000 /* 0x8268 */;
                8347: data_o = 32'h00000000 /* 0x826c */;
                8348: data_o = 32'h00000000 /* 0x8270 */;
                8349: data_o = 32'h00000000 /* 0x8274 */;
                8350: data_o = 32'h00000000 /* 0x8278 */;
                8351: data_o = 32'h00000000 /* 0x827c */;
                8352: data_o = 32'h00000000 /* 0x8280 */;
                8353: data_o = 32'h00000000 /* 0x8284 */;
                8354: data_o = 32'h00000000 /* 0x8288 */;
                8355: data_o = 32'h00000000 /* 0x828c */;
                8356: data_o = 32'h00000000 /* 0x8290 */;
                8357: data_o = 32'h00000000 /* 0x8294 */;
                8358: data_o = 32'h00000000 /* 0x8298 */;
                8359: data_o = 32'h00000000 /* 0x829c */;
                8360: data_o = 32'h00000000 /* 0x82a0 */;
                8361: data_o = 32'h00000000 /* 0x82a4 */;
                8362: data_o = 32'h00000000 /* 0x82a8 */;
                8363: data_o = 32'h00000000 /* 0x82ac */;
                8364: data_o = 32'h00000000 /* 0x82b0 */;
                8365: data_o = 32'h00000000 /* 0x82b4 */;
                8366: data_o = 32'h00000000 /* 0x82b8 */;
                8367: data_o = 32'h00000000 /* 0x82bc */;
                8368: data_o = 32'h00000000 /* 0x82c0 */;
                8369: data_o = 32'h00000000 /* 0x82c4 */;
                8370: data_o = 32'h00000000 /* 0x82c8 */;
                8371: data_o = 32'h00000000 /* 0x82cc */;
                8372: data_o = 32'h00000000 /* 0x82d0 */;
                8373: data_o = 32'h00000000 /* 0x82d4 */;
                8374: data_o = 32'h00000000 /* 0x82d8 */;
                8375: data_o = 32'h00000000 /* 0x82dc */;
                8376: data_o = 32'h00000000 /* 0x82e0 */;
                8377: data_o = 32'h00000000 /* 0x82e4 */;
                8378: data_o = 32'h00000000 /* 0x82e8 */;
                8379: data_o = 32'h00000000 /* 0x82ec */;
                8380: data_o = 32'h00000000 /* 0x82f0 */;
                8381: data_o = 32'h00000000 /* 0x82f4 */;
                8382: data_o = 32'h00000000 /* 0x82f8 */;
                8383: data_o = 32'h00000000 /* 0x82fc */;
                8384: data_o = 32'h00000000 /* 0x8300 */;
                8385: data_o = 32'h00000000 /* 0x8304 */;
                8386: data_o = 32'h00000000 /* 0x8308 */;
                8387: data_o = 32'h00000000 /* 0x830c */;
                8388: data_o = 32'h00000000 /* 0x8310 */;
                8389: data_o = 32'h00000000 /* 0x8314 */;
                8390: data_o = 32'h00000000 /* 0x8318 */;
                8391: data_o = 32'h00000000 /* 0x831c */;
                8392: data_o = 32'h00000000 /* 0x8320 */;
                8393: data_o = 32'h00000000 /* 0x8324 */;
                8394: data_o = 32'h00000000 /* 0x8328 */;
                8395: data_o = 32'h00000000 /* 0x832c */;
                8396: data_o = 32'h00000000 /* 0x8330 */;
                8397: data_o = 32'h00000000 /* 0x8334 */;
                8398: data_o = 32'h00000000 /* 0x8338 */;
                8399: data_o = 32'h00000000 /* 0x833c */;
                8400: data_o = 32'h00000000 /* 0x8340 */;
                8401: data_o = 32'h00000000 /* 0x8344 */;
                8402: data_o = 32'h00000000 /* 0x8348 */;
                8403: data_o = 32'h00000000 /* 0x834c */;
                8404: data_o = 32'h00000000 /* 0x8350 */;
                8405: data_o = 32'h00000000 /* 0x8354 */;
                8406: data_o = 32'h00000000 /* 0x8358 */;
                8407: data_o = 32'h00000000 /* 0x835c */;
                8408: data_o = 32'h00000000 /* 0x8360 */;
                8409: data_o = 32'h00000000 /* 0x8364 */;
                8410: data_o = 32'h00000000 /* 0x8368 */;
                8411: data_o = 32'h00000000 /* 0x836c */;
                8412: data_o = 32'h00000000 /* 0x8370 */;
                8413: data_o = 32'h00000000 /* 0x8374 */;
                8414: data_o = 32'h00000000 /* 0x8378 */;
                8415: data_o = 32'h00000000 /* 0x837c */;
                8416: data_o = 32'h00000000 /* 0x8380 */;
                8417: data_o = 32'h00000000 /* 0x8384 */;
                8418: data_o = 32'h00000000 /* 0x8388 */;
                8419: data_o = 32'h00000000 /* 0x838c */;
                8420: data_o = 32'h00000000 /* 0x8390 */;
                8421: data_o = 32'h00000000 /* 0x8394 */;
                8422: data_o = 32'h00000000 /* 0x8398 */;
                8423: data_o = 32'h00000000 /* 0x839c */;
                8424: data_o = 32'h00000000 /* 0x83a0 */;
                8425: data_o = 32'h00000000 /* 0x83a4 */;
                8426: data_o = 32'h00000000 /* 0x83a8 */;
                8427: data_o = 32'h00000000 /* 0x83ac */;
                8428: data_o = 32'h00000000 /* 0x83b0 */;
                8429: data_o = 32'h00000000 /* 0x83b4 */;
                8430: data_o = 32'h00000000 /* 0x83b8 */;
                8431: data_o = 32'h00000000 /* 0x83bc */;
                8432: data_o = 32'h00000000 /* 0x83c0 */;
                8433: data_o = 32'h00000000 /* 0x83c4 */;
                8434: data_o = 32'h00000000 /* 0x83c8 */;
                8435: data_o = 32'h00000000 /* 0x83cc */;
                8436: data_o = 32'h00000000 /* 0x83d0 */;
                8437: data_o = 32'h00000000 /* 0x83d4 */;
                8438: data_o = 32'h00000000 /* 0x83d8 */;
                8439: data_o = 32'h00000000 /* 0x83dc */;
                8440: data_o = 32'h00000000 /* 0x83e0 */;
                8441: data_o = 32'h00000000 /* 0x83e4 */;
                8442: data_o = 32'h00000000 /* 0x83e8 */;
                8443: data_o = 32'h00000000 /* 0x83ec */;
                8444: data_o = 32'h00000000 /* 0x83f0 */;
                8445: data_o = 32'h00000000 /* 0x83f4 */;
                8446: data_o = 32'h00000000 /* 0x83f8 */;
                8447: data_o = 32'h00000000 /* 0x83fc */;
                8448: data_o = 32'h00000000 /* 0x8400 */;
                8449: data_o = 32'h00000000 /* 0x8404 */;
                8450: data_o = 32'h00000000 /* 0x8408 */;
                8451: data_o = 32'h00000000 /* 0x840c */;
                8452: data_o = 32'h00000000 /* 0x8410 */;
                8453: data_o = 32'h00000000 /* 0x8414 */;
                8454: data_o = 32'h00000000 /* 0x8418 */;
                8455: data_o = 32'h00000000 /* 0x841c */;
                8456: data_o = 32'h00000000 /* 0x8420 */;
                8457: data_o = 32'h00000000 /* 0x8424 */;
                8458: data_o = 32'h00000000 /* 0x8428 */;
                8459: data_o = 32'h00000000 /* 0x842c */;
                8460: data_o = 32'h00000000 /* 0x8430 */;
                8461: data_o = 32'h00000000 /* 0x8434 */;
                8462: data_o = 32'h00000000 /* 0x8438 */;
                8463: data_o = 32'h00000000 /* 0x843c */;
                8464: data_o = 32'h00000000 /* 0x8440 */;
                8465: data_o = 32'h00000000 /* 0x8444 */;
                8466: data_o = 32'h00000000 /* 0x8448 */;
                8467: data_o = 32'h00000000 /* 0x844c */;
                8468: data_o = 32'h00000000 /* 0x8450 */;
                8469: data_o = 32'h00000000 /* 0x8454 */;
                8470: data_o = 32'h00000000 /* 0x8458 */;
                8471: data_o = 32'h00000000 /* 0x845c */;
                8472: data_o = 32'h00000000 /* 0x8460 */;
                8473: data_o = 32'h00000000 /* 0x8464 */;
                8474: data_o = 32'h00000000 /* 0x8468 */;
                8475: data_o = 32'h00000000 /* 0x846c */;
                8476: data_o = 32'h00000000 /* 0x8470 */;
                8477: data_o = 32'h00000000 /* 0x8474 */;
                8478: data_o = 32'h00000000 /* 0x8478 */;
                8479: data_o = 32'h00000000 /* 0x847c */;
                8480: data_o = 32'h00000000 /* 0x8480 */;
                8481: data_o = 32'h00000000 /* 0x8484 */;
                8482: data_o = 32'h00000000 /* 0x8488 */;
                8483: data_o = 32'h00000000 /* 0x848c */;
                8484: data_o = 32'h00000000 /* 0x8490 */;
                8485: data_o = 32'h00000000 /* 0x8494 */;
                8486: data_o = 32'h00000000 /* 0x8498 */;
                8487: data_o = 32'h00000000 /* 0x849c */;
                8488: data_o = 32'h00000000 /* 0x84a0 */;
                8489: data_o = 32'h00000000 /* 0x84a4 */;
                8490: data_o = 32'h00000000 /* 0x84a8 */;
                8491: data_o = 32'h00000000 /* 0x84ac */;
                8492: data_o = 32'h00000000 /* 0x84b0 */;
                8493: data_o = 32'h00000000 /* 0x84b4 */;
                8494: data_o = 32'h00000000 /* 0x84b8 */;
                8495: data_o = 32'h00000000 /* 0x84bc */;
                8496: data_o = 32'h00000000 /* 0x84c0 */;
                8497: data_o = 32'h00000000 /* 0x84c4 */;
                8498: data_o = 32'h00000000 /* 0x84c8 */;
                8499: data_o = 32'h00000000 /* 0x84cc */;
                8500: data_o = 32'h00000000 /* 0x84d0 */;
                8501: data_o = 32'h00000000 /* 0x84d4 */;
                8502: data_o = 32'h00000000 /* 0x84d8 */;
                8503: data_o = 32'h00000000 /* 0x84dc */;
                8504: data_o = 32'h00000000 /* 0x84e0 */;
                8505: data_o = 32'h00000000 /* 0x84e4 */;
                8506: data_o = 32'h00000000 /* 0x84e8 */;
                8507: data_o = 32'h00000000 /* 0x84ec */;
                8508: data_o = 32'h00000000 /* 0x84f0 */;
                8509: data_o = 32'h00000000 /* 0x84f4 */;
                8510: data_o = 32'h00000000 /* 0x84f8 */;
                8511: data_o = 32'h00000000 /* 0x84fc */;
                8512: data_o = 32'h00000000 /* 0x8500 */;
                8513: data_o = 32'h00000000 /* 0x8504 */;
                8514: data_o = 32'h00000000 /* 0x8508 */;
                8515: data_o = 32'h00000000 /* 0x850c */;
                8516: data_o = 32'h00000000 /* 0x8510 */;
                8517: data_o = 32'h00000000 /* 0x8514 */;
                8518: data_o = 32'h00000000 /* 0x8518 */;
                8519: data_o = 32'h00000000 /* 0x851c */;
                8520: data_o = 32'h00000000 /* 0x8520 */;
                8521: data_o = 32'h00000000 /* 0x8524 */;
                8522: data_o = 32'h00000000 /* 0x8528 */;
                8523: data_o = 32'h00000000 /* 0x852c */;
                8524: data_o = 32'h00000000 /* 0x8530 */;
                8525: data_o = 32'h00000000 /* 0x8534 */;
                8526: data_o = 32'h00000000 /* 0x8538 */;
                8527: data_o = 32'h00000000 /* 0x853c */;
                8528: data_o = 32'h00000000 /* 0x8540 */;
                8529: data_o = 32'h00000000 /* 0x8544 */;
                8530: data_o = 32'h00000000 /* 0x8548 */;
                8531: data_o = 32'h00000000 /* 0x854c */;
                8532: data_o = 32'h00000000 /* 0x8550 */;
                8533: data_o = 32'h00000000 /* 0x8554 */;
                8534: data_o = 32'h00000000 /* 0x8558 */;
                8535: data_o = 32'h00000000 /* 0x855c */;
                8536: data_o = 32'h00000000 /* 0x8560 */;
                8537: data_o = 32'h00000000 /* 0x8564 */;
                8538: data_o = 32'h00000000 /* 0x8568 */;
                8539: data_o = 32'h00000000 /* 0x856c */;
                8540: data_o = 32'h00000000 /* 0x8570 */;
                8541: data_o = 32'h00000000 /* 0x8574 */;
                8542: data_o = 32'h00000000 /* 0x8578 */;
                8543: data_o = 32'h00000000 /* 0x857c */;
                8544: data_o = 32'h00000000 /* 0x8580 */;
                8545: data_o = 32'h00000000 /* 0x8584 */;
                8546: data_o = 32'h00000000 /* 0x8588 */;
                8547: data_o = 32'h00000000 /* 0x858c */;
                8548: data_o = 32'h00000000 /* 0x8590 */;
                8549: data_o = 32'h00000000 /* 0x8594 */;
                8550: data_o = 32'h00000000 /* 0x8598 */;
                8551: data_o = 32'h00000000 /* 0x859c */;
                8552: data_o = 32'h00000000 /* 0x85a0 */;
                8553: data_o = 32'h00000000 /* 0x85a4 */;
                8554: data_o = 32'h00000000 /* 0x85a8 */;
                8555: data_o = 32'h00000000 /* 0x85ac */;
                8556: data_o = 32'h00000000 /* 0x85b0 */;
                8557: data_o = 32'h00000000 /* 0x85b4 */;
                8558: data_o = 32'h00000000 /* 0x85b8 */;
                8559: data_o = 32'h00000000 /* 0x85bc */;
                8560: data_o = 32'h00000000 /* 0x85c0 */;
                8561: data_o = 32'h00000000 /* 0x85c4 */;
                8562: data_o = 32'h00000000 /* 0x85c8 */;
                8563: data_o = 32'h00000000 /* 0x85cc */;
                8564: data_o = 32'h00000000 /* 0x85d0 */;
                8565: data_o = 32'h00000000 /* 0x85d4 */;
                8566: data_o = 32'h00000000 /* 0x85d8 */;
                8567: data_o = 32'h00000000 /* 0x85dc */;
                8568: data_o = 32'h00000000 /* 0x85e0 */;
                8569: data_o = 32'h00000000 /* 0x85e4 */;
                8570: data_o = 32'h00000000 /* 0x85e8 */;
                8571: data_o = 32'h00000000 /* 0x85ec */;
                8572: data_o = 32'h00000000 /* 0x85f0 */;
                8573: data_o = 32'h00000000 /* 0x85f4 */;
                8574: data_o = 32'h00000000 /* 0x85f8 */;
                8575: data_o = 32'h00000000 /* 0x85fc */;
                8576: data_o = 32'h00000000 /* 0x8600 */;
                8577: data_o = 32'h00000000 /* 0x8604 */;
                8578: data_o = 32'h00000000 /* 0x8608 */;
                8579: data_o = 32'h00000000 /* 0x860c */;
                8580: data_o = 32'h00000000 /* 0x8610 */;
                8581: data_o = 32'h00000000 /* 0x8614 */;
                8582: data_o = 32'h00000000 /* 0x8618 */;
                8583: data_o = 32'h00000000 /* 0x861c */;
                8584: data_o = 32'h00000000 /* 0x8620 */;
                8585: data_o = 32'h00000000 /* 0x8624 */;
                8586: data_o = 32'h00000000 /* 0x8628 */;
                8587: data_o = 32'h00000000 /* 0x862c */;
                8588: data_o = 32'h00000000 /* 0x8630 */;
                8589: data_o = 32'h00000000 /* 0x8634 */;
                8590: data_o = 32'h00000000 /* 0x8638 */;
                8591: data_o = 32'h00000000 /* 0x863c */;
                8592: data_o = 32'h00000000 /* 0x8640 */;
                8593: data_o = 32'h00000000 /* 0x8644 */;
                8594: data_o = 32'h00000000 /* 0x8648 */;
                8595: data_o = 32'h00000000 /* 0x864c */;
                8596: data_o = 32'h00000000 /* 0x8650 */;
                8597: data_o = 32'h00000000 /* 0x8654 */;
                8598: data_o = 32'h00000000 /* 0x8658 */;
                8599: data_o = 32'h00000000 /* 0x865c */;
                8600: data_o = 32'h00000000 /* 0x8660 */;
                8601: data_o = 32'h00000000 /* 0x8664 */;
                8602: data_o = 32'h00000000 /* 0x8668 */;
                8603: data_o = 32'h00000000 /* 0x866c */;
                8604: data_o = 32'h00000000 /* 0x8670 */;
                8605: data_o = 32'h00000000 /* 0x8674 */;
                8606: data_o = 32'h00000000 /* 0x8678 */;
                8607: data_o = 32'h00000000 /* 0x867c */;
                8608: data_o = 32'h00000000 /* 0x8680 */;
                8609: data_o = 32'h00000000 /* 0x8684 */;
                8610: data_o = 32'h00000000 /* 0x8688 */;
                8611: data_o = 32'h00000000 /* 0x868c */;
                8612: data_o = 32'h00000000 /* 0x8690 */;
                8613: data_o = 32'h00000000 /* 0x8694 */;
                8614: data_o = 32'h00000000 /* 0x8698 */;
                8615: data_o = 32'h00000000 /* 0x869c */;
                8616: data_o = 32'h00000000 /* 0x86a0 */;
                8617: data_o = 32'h00000000 /* 0x86a4 */;
                8618: data_o = 32'h00000000 /* 0x86a8 */;
                8619: data_o = 32'h00000000 /* 0x86ac */;
                8620: data_o = 32'h00000000 /* 0x86b0 */;
                8621: data_o = 32'h00000000 /* 0x86b4 */;
                8622: data_o = 32'h00000000 /* 0x86b8 */;
                8623: data_o = 32'h00000000 /* 0x86bc */;
                8624: data_o = 32'h00000000 /* 0x86c0 */;
                8625: data_o = 32'h00000000 /* 0x86c4 */;
                8626: data_o = 32'h00000000 /* 0x86c8 */;
                8627: data_o = 32'h00000000 /* 0x86cc */;
                8628: data_o = 32'h00000000 /* 0x86d0 */;
                8629: data_o = 32'h00000000 /* 0x86d4 */;
                8630: data_o = 32'h00000000 /* 0x86d8 */;
                8631: data_o = 32'h00000000 /* 0x86dc */;
                8632: data_o = 32'h00000000 /* 0x86e0 */;
                8633: data_o = 32'h00000000 /* 0x86e4 */;
                8634: data_o = 32'h00000000 /* 0x86e8 */;
                8635: data_o = 32'h00000000 /* 0x86ec */;
                8636: data_o = 32'h00000000 /* 0x86f0 */;
                8637: data_o = 32'h00000000 /* 0x86f4 */;
                8638: data_o = 32'h00000000 /* 0x86f8 */;
                8639: data_o = 32'h00000000 /* 0x86fc */;
                8640: data_o = 32'h00000000 /* 0x8700 */;
                8641: data_o = 32'h00000000 /* 0x8704 */;
                8642: data_o = 32'h00000000 /* 0x8708 */;
                8643: data_o = 32'h00000000 /* 0x870c */;
                8644: data_o = 32'h00000000 /* 0x8710 */;
                8645: data_o = 32'h00000000 /* 0x8714 */;
                8646: data_o = 32'h00000000 /* 0x8718 */;
                8647: data_o = 32'h00000000 /* 0x871c */;
                8648: data_o = 32'h00000000 /* 0x8720 */;
                8649: data_o = 32'h00000000 /* 0x8724 */;
                8650: data_o = 32'h00000000 /* 0x8728 */;
                8651: data_o = 32'h00000000 /* 0x872c */;
                8652: data_o = 32'h00000000 /* 0x8730 */;
                8653: data_o = 32'h00000000 /* 0x8734 */;
                8654: data_o = 32'h00000000 /* 0x8738 */;
                8655: data_o = 32'h00000000 /* 0x873c */;
                8656: data_o = 32'h00000000 /* 0x8740 */;
                8657: data_o = 32'h00000000 /* 0x8744 */;
                8658: data_o = 32'h00000000 /* 0x8748 */;
                8659: data_o = 32'h00000000 /* 0x874c */;
                8660: data_o = 32'h00000000 /* 0x8750 */;
                8661: data_o = 32'h00000000 /* 0x8754 */;
                8662: data_o = 32'h00000000 /* 0x8758 */;
                8663: data_o = 32'h00000000 /* 0x875c */;
                8664: data_o = 32'h00000000 /* 0x8760 */;
                8665: data_o = 32'h00000000 /* 0x8764 */;
                8666: data_o = 32'h00000000 /* 0x8768 */;
                8667: data_o = 32'h00000000 /* 0x876c */;
                8668: data_o = 32'h00000000 /* 0x8770 */;
                8669: data_o = 32'h00000000 /* 0x8774 */;
                8670: data_o = 32'h00000000 /* 0x8778 */;
                8671: data_o = 32'h00000000 /* 0x877c */;
                8672: data_o = 32'h00000000 /* 0x8780 */;
                8673: data_o = 32'h00000000 /* 0x8784 */;
                8674: data_o = 32'h00000000 /* 0x8788 */;
                8675: data_o = 32'h00000000 /* 0x878c */;
                8676: data_o = 32'h00000000 /* 0x8790 */;
                8677: data_o = 32'h00000000 /* 0x8794 */;
                8678: data_o = 32'h00000000 /* 0x8798 */;
                8679: data_o = 32'h00000000 /* 0x879c */;
                8680: data_o = 32'h00000000 /* 0x87a0 */;
                8681: data_o = 32'h00000000 /* 0x87a4 */;
                8682: data_o = 32'h00000000 /* 0x87a8 */;
                8683: data_o = 32'h00000000 /* 0x87ac */;
                8684: data_o = 32'h00000000 /* 0x87b0 */;
                8685: data_o = 32'h00000000 /* 0x87b4 */;
                8686: data_o = 32'h00000000 /* 0x87b8 */;
                8687: data_o = 32'h00000000 /* 0x87bc */;
                8688: data_o = 32'h00000000 /* 0x87c0 */;
                8689: data_o = 32'h00000000 /* 0x87c4 */;
                8690: data_o = 32'h00000000 /* 0x87c8 */;
                8691: data_o = 32'h00000000 /* 0x87cc */;
                8692: data_o = 32'h00000000 /* 0x87d0 */;
                8693: data_o = 32'h00000000 /* 0x87d4 */;
                8694: data_o = 32'h00000000 /* 0x87d8 */;
                8695: data_o = 32'h00000000 /* 0x87dc */;
                8696: data_o = 32'h00000000 /* 0x87e0 */;
                8697: data_o = 32'h00000000 /* 0x87e4 */;
                8698: data_o = 32'h00000000 /* 0x87e8 */;
                8699: data_o = 32'h00000000 /* 0x87ec */;
                8700: data_o = 32'h00000000 /* 0x87f0 */;
                8701: data_o = 32'h00000000 /* 0x87f4 */;
                8702: data_o = 32'h00000000 /* 0x87f8 */;
                8703: data_o = 32'h00000000 /* 0x87fc */;
                8704: data_o = 32'h00000000 /* 0x8800 */;
                8705: data_o = 32'h00000000 /* 0x8804 */;
                8706: data_o = 32'h00000000 /* 0x8808 */;
                8707: data_o = 32'h00000000 /* 0x880c */;
                8708: data_o = 32'h00000000 /* 0x8810 */;
                8709: data_o = 32'h00000000 /* 0x8814 */;
                8710: data_o = 32'h00000000 /* 0x8818 */;
                8711: data_o = 32'h00000000 /* 0x881c */;
                8712: data_o = 32'h00000000 /* 0x8820 */;
                8713: data_o = 32'h00000000 /* 0x8824 */;
                8714: data_o = 32'h00000000 /* 0x8828 */;
                8715: data_o = 32'h00000000 /* 0x882c */;
                8716: data_o = 32'h00000000 /* 0x8830 */;
                8717: data_o = 32'h00000000 /* 0x8834 */;
                8718: data_o = 32'h00000000 /* 0x8838 */;
                8719: data_o = 32'h00000000 /* 0x883c */;
                8720: data_o = 32'h00000000 /* 0x8840 */;
                8721: data_o = 32'h00000000 /* 0x8844 */;
                8722: data_o = 32'h00000000 /* 0x8848 */;
                8723: data_o = 32'h00000000 /* 0x884c */;
                8724: data_o = 32'h00000000 /* 0x8850 */;
                8725: data_o = 32'h00000000 /* 0x8854 */;
                8726: data_o = 32'h00000000 /* 0x8858 */;
                8727: data_o = 32'h00000000 /* 0x885c */;
                8728: data_o = 32'h00000000 /* 0x8860 */;
                8729: data_o = 32'h00000000 /* 0x8864 */;
                8730: data_o = 32'h00000000 /* 0x8868 */;
                8731: data_o = 32'h00000000 /* 0x886c */;
                8732: data_o = 32'h00000000 /* 0x8870 */;
                8733: data_o = 32'h00000000 /* 0x8874 */;
                8734: data_o = 32'h00000000 /* 0x8878 */;
                8735: data_o = 32'h00000000 /* 0x887c */;
                8736: data_o = 32'h00000000 /* 0x8880 */;
                8737: data_o = 32'h00000000 /* 0x8884 */;
                8738: data_o = 32'h00000000 /* 0x8888 */;
                8739: data_o = 32'h00000000 /* 0x888c */;
                8740: data_o = 32'h00000000 /* 0x8890 */;
                8741: data_o = 32'h00000000 /* 0x8894 */;
                8742: data_o = 32'h00000000 /* 0x8898 */;
                8743: data_o = 32'h00000000 /* 0x889c */;
                8744: data_o = 32'h00000000 /* 0x88a0 */;
                8745: data_o = 32'h00000000 /* 0x88a4 */;
                8746: data_o = 32'h00000000 /* 0x88a8 */;
                8747: data_o = 32'h00000000 /* 0x88ac */;
                8748: data_o = 32'h00000000 /* 0x88b0 */;
                8749: data_o = 32'h00000000 /* 0x88b4 */;
                8750: data_o = 32'h00000000 /* 0x88b8 */;
                8751: data_o = 32'h00000000 /* 0x88bc */;
                8752: data_o = 32'h00000000 /* 0x88c0 */;
                8753: data_o = 32'h00000000 /* 0x88c4 */;
                8754: data_o = 32'h00000000 /* 0x88c8 */;
                8755: data_o = 32'h00000000 /* 0x88cc */;
                8756: data_o = 32'h00000000 /* 0x88d0 */;
                8757: data_o = 32'h00000000 /* 0x88d4 */;
                8758: data_o = 32'h00000000 /* 0x88d8 */;
                8759: data_o = 32'h00000000 /* 0x88dc */;
                8760: data_o = 32'h00000000 /* 0x88e0 */;
                8761: data_o = 32'h00000000 /* 0x88e4 */;
                8762: data_o = 32'h00000000 /* 0x88e8 */;
                8763: data_o = 32'h00000000 /* 0x88ec */;
                8764: data_o = 32'h00000000 /* 0x88f0 */;
                8765: data_o = 32'h00000000 /* 0x88f4 */;
                8766: data_o = 32'h00000000 /* 0x88f8 */;
                8767: data_o = 32'h00000000 /* 0x88fc */;
                8768: data_o = 32'h00000000 /* 0x8900 */;
                8769: data_o = 32'h00000000 /* 0x8904 */;
                8770: data_o = 32'h00000000 /* 0x8908 */;
                8771: data_o = 32'h00000000 /* 0x890c */;
                8772: data_o = 32'h00000000 /* 0x8910 */;
                8773: data_o = 32'h00000000 /* 0x8914 */;
                8774: data_o = 32'h00000000 /* 0x8918 */;
                8775: data_o = 32'h00000000 /* 0x891c */;
                8776: data_o = 32'h00000000 /* 0x8920 */;
                8777: data_o = 32'h00000000 /* 0x8924 */;
                8778: data_o = 32'h00000000 /* 0x8928 */;
                8779: data_o = 32'h00000000 /* 0x892c */;
                8780: data_o = 32'h00000000 /* 0x8930 */;
                8781: data_o = 32'h00000000 /* 0x8934 */;
                8782: data_o = 32'h00000000 /* 0x8938 */;
                8783: data_o = 32'h00000000 /* 0x893c */;
                8784: data_o = 32'h00000000 /* 0x8940 */;
                8785: data_o = 32'h00000000 /* 0x8944 */;
                8786: data_o = 32'h00000000 /* 0x8948 */;
                8787: data_o = 32'h00000000 /* 0x894c */;
                8788: data_o = 32'h00000000 /* 0x8950 */;
                8789: data_o = 32'h00000000 /* 0x8954 */;
                8790: data_o = 32'h00000000 /* 0x8958 */;
                8791: data_o = 32'h00000000 /* 0x895c */;
                8792: data_o = 32'h00000000 /* 0x8960 */;
                8793: data_o = 32'h00000000 /* 0x8964 */;
                8794: data_o = 32'h00000000 /* 0x8968 */;
                8795: data_o = 32'h00000000 /* 0x896c */;
                8796: data_o = 32'h00000000 /* 0x8970 */;
                8797: data_o = 32'h00000000 /* 0x8974 */;
                8798: data_o = 32'h00000000 /* 0x8978 */;
                8799: data_o = 32'h00000000 /* 0x897c */;
                8800: data_o = 32'h00000000 /* 0x8980 */;
                8801: data_o = 32'h00000000 /* 0x8984 */;
                8802: data_o = 32'h00000000 /* 0x8988 */;
                8803: data_o = 32'h00000000 /* 0x898c */;
                8804: data_o = 32'h00000000 /* 0x8990 */;
                8805: data_o = 32'h00000000 /* 0x8994 */;
                8806: data_o = 32'h00000000 /* 0x8998 */;
                8807: data_o = 32'h00000000 /* 0x899c */;
                8808: data_o = 32'h00000000 /* 0x89a0 */;
                8809: data_o = 32'h00000000 /* 0x89a4 */;
                8810: data_o = 32'h00000000 /* 0x89a8 */;
                8811: data_o = 32'h00000000 /* 0x89ac */;
                8812: data_o = 32'h00000000 /* 0x89b0 */;
                8813: data_o = 32'h00000000 /* 0x89b4 */;
                8814: data_o = 32'h00000000 /* 0x89b8 */;
                8815: data_o = 32'h00000000 /* 0x89bc */;
                8816: data_o = 32'h00000000 /* 0x89c0 */;
                8817: data_o = 32'h00000000 /* 0x89c4 */;
                8818: data_o = 32'h00000000 /* 0x89c8 */;
                8819: data_o = 32'h00000000 /* 0x89cc */;
                8820: data_o = 32'h00000000 /* 0x89d0 */;
                8821: data_o = 32'h00000000 /* 0x89d4 */;
                8822: data_o = 32'h00000000 /* 0x89d8 */;
                8823: data_o = 32'h00000000 /* 0x89dc */;
                8824: data_o = 32'h00000000 /* 0x89e0 */;
                8825: data_o = 32'h00000000 /* 0x89e4 */;
                8826: data_o = 32'h00000000 /* 0x89e8 */;
                8827: data_o = 32'h00000000 /* 0x89ec */;
                8828: data_o = 32'h00000000 /* 0x89f0 */;
                8829: data_o = 32'h00000000 /* 0x89f4 */;
                8830: data_o = 32'h00000000 /* 0x89f8 */;
                8831: data_o = 32'h00000000 /* 0x89fc */;
                8832: data_o = 32'h00000000 /* 0x8a00 */;
                8833: data_o = 32'h00000000 /* 0x8a04 */;
                8834: data_o = 32'h00000000 /* 0x8a08 */;
                8835: data_o = 32'h00000000 /* 0x8a0c */;
                8836: data_o = 32'h00000000 /* 0x8a10 */;
                8837: data_o = 32'h00000000 /* 0x8a14 */;
                8838: data_o = 32'h00000000 /* 0x8a18 */;
                8839: data_o = 32'h00000000 /* 0x8a1c */;
                8840: data_o = 32'h00000000 /* 0x8a20 */;
                8841: data_o = 32'h00000000 /* 0x8a24 */;
                8842: data_o = 32'h00000000 /* 0x8a28 */;
                8843: data_o = 32'h00000000 /* 0x8a2c */;
                8844: data_o = 32'h00000000 /* 0x8a30 */;
                8845: data_o = 32'h00000000 /* 0x8a34 */;
                8846: data_o = 32'h00000000 /* 0x8a38 */;
                8847: data_o = 32'h00000000 /* 0x8a3c */;
                8848: data_o = 32'h00000000 /* 0x8a40 */;
                8849: data_o = 32'h00000000 /* 0x8a44 */;
                8850: data_o = 32'h00000000 /* 0x8a48 */;
                8851: data_o = 32'h00000000 /* 0x8a4c */;
                8852: data_o = 32'h00000000 /* 0x8a50 */;
                8853: data_o = 32'h00000000 /* 0x8a54 */;
                8854: data_o = 32'h00000000 /* 0x8a58 */;
                8855: data_o = 32'h00000000 /* 0x8a5c */;
                8856: data_o = 32'h00000000 /* 0x8a60 */;
                8857: data_o = 32'h00000000 /* 0x8a64 */;
                8858: data_o = 32'h00000000 /* 0x8a68 */;
                8859: data_o = 32'h00000000 /* 0x8a6c */;
                8860: data_o = 32'h00000000 /* 0x8a70 */;
                8861: data_o = 32'h00000000 /* 0x8a74 */;
                8862: data_o = 32'h00000000 /* 0x8a78 */;
                8863: data_o = 32'h00000000 /* 0x8a7c */;
                8864: data_o = 32'h00000000 /* 0x8a80 */;
                8865: data_o = 32'h00000000 /* 0x8a84 */;
                8866: data_o = 32'h00000000 /* 0x8a88 */;
                8867: data_o = 32'h00000000 /* 0x8a8c */;
                8868: data_o = 32'h00000000 /* 0x8a90 */;
                8869: data_o = 32'h00000000 /* 0x8a94 */;
                8870: data_o = 32'h00000000 /* 0x8a98 */;
                8871: data_o = 32'h00000000 /* 0x8a9c */;
                8872: data_o = 32'h00000000 /* 0x8aa0 */;
                8873: data_o = 32'h00000000 /* 0x8aa4 */;
                8874: data_o = 32'h00000000 /* 0x8aa8 */;
                8875: data_o = 32'h00000000 /* 0x8aac */;
                8876: data_o = 32'h00000000 /* 0x8ab0 */;
                8877: data_o = 32'h00000000 /* 0x8ab4 */;
                8878: data_o = 32'h00000000 /* 0x8ab8 */;
                8879: data_o = 32'h00000000 /* 0x8abc */;
                8880: data_o = 32'h00000000 /* 0x8ac0 */;
                8881: data_o = 32'h00000000 /* 0x8ac4 */;
                8882: data_o = 32'h00000000 /* 0x8ac8 */;
                8883: data_o = 32'h00000000 /* 0x8acc */;
                8884: data_o = 32'h00000000 /* 0x8ad0 */;
                8885: data_o = 32'h00000000 /* 0x8ad4 */;
                8886: data_o = 32'h00000000 /* 0x8ad8 */;
                8887: data_o = 32'h00000000 /* 0x8adc */;
                8888: data_o = 32'h00000000 /* 0x8ae0 */;
                8889: data_o = 32'h00000000 /* 0x8ae4 */;
                8890: data_o = 32'h00000000 /* 0x8ae8 */;
                8891: data_o = 32'h00000000 /* 0x8aec */;
                8892: data_o = 32'h00000000 /* 0x8af0 */;
                8893: data_o = 32'h00000000 /* 0x8af4 */;
                8894: data_o = 32'h00000000 /* 0x8af8 */;
                8895: data_o = 32'h00000000 /* 0x8afc */;
                8896: data_o = 32'h00000000 /* 0x8b00 */;
                8897: data_o = 32'h00000000 /* 0x8b04 */;
                8898: data_o = 32'h00000000 /* 0x8b08 */;
                8899: data_o = 32'h00000000 /* 0x8b0c */;
                8900: data_o = 32'h00000000 /* 0x8b10 */;
                8901: data_o = 32'h00000000 /* 0x8b14 */;
                8902: data_o = 32'h00000000 /* 0x8b18 */;
                8903: data_o = 32'h00000000 /* 0x8b1c */;
                8904: data_o = 32'h00000000 /* 0x8b20 */;
                8905: data_o = 32'h00000000 /* 0x8b24 */;
                8906: data_o = 32'h00000000 /* 0x8b28 */;
                8907: data_o = 32'h00000000 /* 0x8b2c */;
                8908: data_o = 32'h00000000 /* 0x8b30 */;
                8909: data_o = 32'h00000000 /* 0x8b34 */;
                8910: data_o = 32'h00000000 /* 0x8b38 */;
                8911: data_o = 32'h00000000 /* 0x8b3c */;
                8912: data_o = 32'h00000000 /* 0x8b40 */;
                8913: data_o = 32'h00000000 /* 0x8b44 */;
                8914: data_o = 32'h00000000 /* 0x8b48 */;
                8915: data_o = 32'h00000000 /* 0x8b4c */;
                8916: data_o = 32'h00000000 /* 0x8b50 */;
                8917: data_o = 32'h00000000 /* 0x8b54 */;
                8918: data_o = 32'h00000000 /* 0x8b58 */;
                8919: data_o = 32'h00000000 /* 0x8b5c */;
                8920: data_o = 32'h00000000 /* 0x8b60 */;
                8921: data_o = 32'h00000000 /* 0x8b64 */;
                8922: data_o = 32'h00000000 /* 0x8b68 */;
                8923: data_o = 32'h00000000 /* 0x8b6c */;
                8924: data_o = 32'h00000000 /* 0x8b70 */;
                8925: data_o = 32'h00000000 /* 0x8b74 */;
                8926: data_o = 32'h00000000 /* 0x8b78 */;
                8927: data_o = 32'h00000000 /* 0x8b7c */;
                8928: data_o = 32'h00000000 /* 0x8b80 */;
                8929: data_o = 32'h00000000 /* 0x8b84 */;
                8930: data_o = 32'h00000000 /* 0x8b88 */;
                8931: data_o = 32'h00000000 /* 0x8b8c */;
                8932: data_o = 32'h00000000 /* 0x8b90 */;
                8933: data_o = 32'h00000000 /* 0x8b94 */;
                8934: data_o = 32'h00000000 /* 0x8b98 */;
                8935: data_o = 32'h00000000 /* 0x8b9c */;
                8936: data_o = 32'h00000000 /* 0x8ba0 */;
                8937: data_o = 32'h00000000 /* 0x8ba4 */;
                8938: data_o = 32'h00000000 /* 0x8ba8 */;
                8939: data_o = 32'h00000000 /* 0x8bac */;
                8940: data_o = 32'h00000000 /* 0x8bb0 */;
                8941: data_o = 32'h00000000 /* 0x8bb4 */;
                8942: data_o = 32'h00000000 /* 0x8bb8 */;
                8943: data_o = 32'h00000000 /* 0x8bbc */;
                8944: data_o = 32'h00000000 /* 0x8bc0 */;
                8945: data_o = 32'h00000000 /* 0x8bc4 */;
                8946: data_o = 32'h00000000 /* 0x8bc8 */;
                8947: data_o = 32'h00000000 /* 0x8bcc */;
                8948: data_o = 32'h00000000 /* 0x8bd0 */;
                8949: data_o = 32'h00000000 /* 0x8bd4 */;
                8950: data_o = 32'h00000000 /* 0x8bd8 */;
                8951: data_o = 32'h00000000 /* 0x8bdc */;
                8952: data_o = 32'h00000000 /* 0x8be0 */;
                8953: data_o = 32'h00000000 /* 0x8be4 */;
                8954: data_o = 32'h00000000 /* 0x8be8 */;
                8955: data_o = 32'h00000000 /* 0x8bec */;
                8956: data_o = 32'h00000000 /* 0x8bf0 */;
                8957: data_o = 32'h00000000 /* 0x8bf4 */;
                8958: data_o = 32'h00000000 /* 0x8bf8 */;
                8959: data_o = 32'h00000000 /* 0x8bfc */;
                8960: data_o = 32'h00000000 /* 0x8c00 */;
                8961: data_o = 32'h00000000 /* 0x8c04 */;
                8962: data_o = 32'h00000000 /* 0x8c08 */;
                8963: data_o = 32'h00000000 /* 0x8c0c */;
                8964: data_o = 32'h00000000 /* 0x8c10 */;
                8965: data_o = 32'h00000000 /* 0x8c14 */;
                8966: data_o = 32'h00000000 /* 0x8c18 */;
                8967: data_o = 32'h00000000 /* 0x8c1c */;
                8968: data_o = 32'h00000000 /* 0x8c20 */;
                8969: data_o = 32'h00000000 /* 0x8c24 */;
                8970: data_o = 32'h00000000 /* 0x8c28 */;
                8971: data_o = 32'h00000000 /* 0x8c2c */;
                8972: data_o = 32'h00000000 /* 0x8c30 */;
                8973: data_o = 32'h00000000 /* 0x8c34 */;
                8974: data_o = 32'h00000000 /* 0x8c38 */;
                8975: data_o = 32'h00000000 /* 0x8c3c */;
                8976: data_o = 32'h00000000 /* 0x8c40 */;
                8977: data_o = 32'h00000000 /* 0x8c44 */;
                8978: data_o = 32'h00000000 /* 0x8c48 */;
                8979: data_o = 32'h00000000 /* 0x8c4c */;
                8980: data_o = 32'h00000000 /* 0x8c50 */;
                8981: data_o = 32'h00000000 /* 0x8c54 */;
                8982: data_o = 32'h00000000 /* 0x8c58 */;
                8983: data_o = 32'h00000000 /* 0x8c5c */;
                8984: data_o = 32'h00000000 /* 0x8c60 */;
                8985: data_o = 32'h00000000 /* 0x8c64 */;
                8986: data_o = 32'h00000000 /* 0x8c68 */;
                8987: data_o = 32'h00000000 /* 0x8c6c */;
                8988: data_o = 32'h00000000 /* 0x8c70 */;
                8989: data_o = 32'h00000000 /* 0x8c74 */;
                8990: data_o = 32'h00000000 /* 0x8c78 */;
                8991: data_o = 32'h00000000 /* 0x8c7c */;
                8992: data_o = 32'h00000000 /* 0x8c80 */;
                8993: data_o = 32'h00000000 /* 0x8c84 */;
                8994: data_o = 32'h00000000 /* 0x8c88 */;
                8995: data_o = 32'h00000000 /* 0x8c8c */;
                8996: data_o = 32'h00000000 /* 0x8c90 */;
                8997: data_o = 32'h00000000 /* 0x8c94 */;
                8998: data_o = 32'h00000000 /* 0x8c98 */;
                8999: data_o = 32'h00000000 /* 0x8c9c */;
                9000: data_o = 32'h00000000 /* 0x8ca0 */;
                9001: data_o = 32'h00000000 /* 0x8ca4 */;
                9002: data_o = 32'h00000000 /* 0x8ca8 */;
                9003: data_o = 32'h00000000 /* 0x8cac */;
                9004: data_o = 32'h00000000 /* 0x8cb0 */;
                9005: data_o = 32'h00000000 /* 0x8cb4 */;
                9006: data_o = 32'h00000000 /* 0x8cb8 */;
                9007: data_o = 32'h00000000 /* 0x8cbc */;
                9008: data_o = 32'h00000000 /* 0x8cc0 */;
                9009: data_o = 32'h00000000 /* 0x8cc4 */;
                9010: data_o = 32'h00000000 /* 0x8cc8 */;
                9011: data_o = 32'h00000000 /* 0x8ccc */;
                9012: data_o = 32'h00000000 /* 0x8cd0 */;
                9013: data_o = 32'h00000000 /* 0x8cd4 */;
                9014: data_o = 32'h00000000 /* 0x8cd8 */;
                9015: data_o = 32'h00000000 /* 0x8cdc */;
                9016: data_o = 32'h00000000 /* 0x8ce0 */;
                9017: data_o = 32'h00000000 /* 0x8ce4 */;
                9018: data_o = 32'h00000000 /* 0x8ce8 */;
                9019: data_o = 32'h00000000 /* 0x8cec */;
                9020: data_o = 32'h00000000 /* 0x8cf0 */;
                9021: data_o = 32'h00000000 /* 0x8cf4 */;
                9022: data_o = 32'h00000000 /* 0x8cf8 */;
                9023: data_o = 32'h00000000 /* 0x8cfc */;
                9024: data_o = 32'h00000000 /* 0x8d00 */;
                9025: data_o = 32'h00000000 /* 0x8d04 */;
                9026: data_o = 32'h00000000 /* 0x8d08 */;
                9027: data_o = 32'h00000000 /* 0x8d0c */;
                9028: data_o = 32'h00000000 /* 0x8d10 */;
                9029: data_o = 32'h00000000 /* 0x8d14 */;
                9030: data_o = 32'h00000000 /* 0x8d18 */;
                9031: data_o = 32'h00000000 /* 0x8d1c */;
                9032: data_o = 32'h00000000 /* 0x8d20 */;
                9033: data_o = 32'h00000000 /* 0x8d24 */;
                9034: data_o = 32'h00000000 /* 0x8d28 */;
                9035: data_o = 32'h00000000 /* 0x8d2c */;
                9036: data_o = 32'h00000000 /* 0x8d30 */;
                9037: data_o = 32'h00000000 /* 0x8d34 */;
                9038: data_o = 32'h00000000 /* 0x8d38 */;
                9039: data_o = 32'h00000000 /* 0x8d3c */;
                9040: data_o = 32'h00000000 /* 0x8d40 */;
                9041: data_o = 32'h00000000 /* 0x8d44 */;
                9042: data_o = 32'h00000000 /* 0x8d48 */;
                9043: data_o = 32'h00000000 /* 0x8d4c */;
                9044: data_o = 32'h00000000 /* 0x8d50 */;
                9045: data_o = 32'h00000000 /* 0x8d54 */;
                9046: data_o = 32'h00000000 /* 0x8d58 */;
                9047: data_o = 32'h00000000 /* 0x8d5c */;
                9048: data_o = 32'h00000000 /* 0x8d60 */;
                9049: data_o = 32'h00000000 /* 0x8d64 */;
                9050: data_o = 32'h00000000 /* 0x8d68 */;
                9051: data_o = 32'h00000000 /* 0x8d6c */;
                9052: data_o = 32'h00000000 /* 0x8d70 */;
                9053: data_o = 32'h00000000 /* 0x8d74 */;
                9054: data_o = 32'h00000000 /* 0x8d78 */;
                9055: data_o = 32'h00000000 /* 0x8d7c */;
                9056: data_o = 32'h00000000 /* 0x8d80 */;
                9057: data_o = 32'h00000000 /* 0x8d84 */;
                9058: data_o = 32'h00000000 /* 0x8d88 */;
                9059: data_o = 32'h00000000 /* 0x8d8c */;
                9060: data_o = 32'h00000000 /* 0x8d90 */;
                9061: data_o = 32'h00000000 /* 0x8d94 */;
                9062: data_o = 32'h00000000 /* 0x8d98 */;
                9063: data_o = 32'h00000000 /* 0x8d9c */;
                9064: data_o = 32'h00000000 /* 0x8da0 */;
                9065: data_o = 32'h00000000 /* 0x8da4 */;
                9066: data_o = 32'h00000000 /* 0x8da8 */;
                9067: data_o = 32'h00000000 /* 0x8dac */;
                9068: data_o = 32'h00000000 /* 0x8db0 */;
                9069: data_o = 32'h00000000 /* 0x8db4 */;
                9070: data_o = 32'h00000000 /* 0x8db8 */;
                9071: data_o = 32'h00000000 /* 0x8dbc */;
                9072: data_o = 32'h00000000 /* 0x8dc0 */;
                9073: data_o = 32'h00000000 /* 0x8dc4 */;
                9074: data_o = 32'h00000000 /* 0x8dc8 */;
                9075: data_o = 32'h00000000 /* 0x8dcc */;
                9076: data_o = 32'h00000000 /* 0x8dd0 */;
                9077: data_o = 32'h00000000 /* 0x8dd4 */;
                9078: data_o = 32'h00000000 /* 0x8dd8 */;
                9079: data_o = 32'h00000000 /* 0x8ddc */;
                9080: data_o = 32'h00000000 /* 0x8de0 */;
                9081: data_o = 32'h00000000 /* 0x8de4 */;
                9082: data_o = 32'h00000000 /* 0x8de8 */;
                9083: data_o = 32'h00000000 /* 0x8dec */;
                9084: data_o = 32'h00000000 /* 0x8df0 */;
                9085: data_o = 32'h00000000 /* 0x8df4 */;
                9086: data_o = 32'h00000000 /* 0x8df8 */;
                9087: data_o = 32'h00000000 /* 0x8dfc */;
                9088: data_o = 32'h00000000 /* 0x8e00 */;
                9089: data_o = 32'h00000000 /* 0x8e04 */;
                9090: data_o = 32'h00000000 /* 0x8e08 */;
                9091: data_o = 32'h00000000 /* 0x8e0c */;
                9092: data_o = 32'h00000000 /* 0x8e10 */;
                9093: data_o = 32'h00000000 /* 0x8e14 */;
                9094: data_o = 32'h00000000 /* 0x8e18 */;
                9095: data_o = 32'h00000000 /* 0x8e1c */;
                9096: data_o = 32'h00000000 /* 0x8e20 */;
                9097: data_o = 32'h00000000 /* 0x8e24 */;
                9098: data_o = 32'h00000000 /* 0x8e28 */;
                9099: data_o = 32'h00000000 /* 0x8e2c */;
                9100: data_o = 32'h00000000 /* 0x8e30 */;
                9101: data_o = 32'h00000000 /* 0x8e34 */;
                9102: data_o = 32'h00000000 /* 0x8e38 */;
                9103: data_o = 32'h00000000 /* 0x8e3c */;
                9104: data_o = 32'h00000000 /* 0x8e40 */;
                9105: data_o = 32'h00000000 /* 0x8e44 */;
                9106: data_o = 32'h00000000 /* 0x8e48 */;
                9107: data_o = 32'h00000000 /* 0x8e4c */;
                9108: data_o = 32'h00000000 /* 0x8e50 */;
                9109: data_o = 32'h00000000 /* 0x8e54 */;
                9110: data_o = 32'h00000000 /* 0x8e58 */;
                9111: data_o = 32'h00000000 /* 0x8e5c */;
                9112: data_o = 32'h00000000 /* 0x8e60 */;
                9113: data_o = 32'h00000000 /* 0x8e64 */;
                9114: data_o = 32'h00000000 /* 0x8e68 */;
                9115: data_o = 32'h00000000 /* 0x8e6c */;
                9116: data_o = 32'h00000000 /* 0x8e70 */;
                9117: data_o = 32'h00000000 /* 0x8e74 */;
                9118: data_o = 32'h00000000 /* 0x8e78 */;
                9119: data_o = 32'h00000000 /* 0x8e7c */;
                9120: data_o = 32'h00000000 /* 0x8e80 */;
                9121: data_o = 32'h00000000 /* 0x8e84 */;
                9122: data_o = 32'h00000000 /* 0x8e88 */;
                9123: data_o = 32'h00000000 /* 0x8e8c */;
                9124: data_o = 32'h00000000 /* 0x8e90 */;
                9125: data_o = 32'h00000000 /* 0x8e94 */;
                9126: data_o = 32'h00000000 /* 0x8e98 */;
                9127: data_o = 32'h00000000 /* 0x8e9c */;
                9128: data_o = 32'h00000000 /* 0x8ea0 */;
                9129: data_o = 32'h00000000 /* 0x8ea4 */;
                9130: data_o = 32'h00000000 /* 0x8ea8 */;
                9131: data_o = 32'h00000000 /* 0x8eac */;
                9132: data_o = 32'h00000000 /* 0x8eb0 */;
                9133: data_o = 32'h00000000 /* 0x8eb4 */;
                9134: data_o = 32'h00000000 /* 0x8eb8 */;
                9135: data_o = 32'h00000000 /* 0x8ebc */;
                9136: data_o = 32'h00000000 /* 0x8ec0 */;
                9137: data_o = 32'h00000000 /* 0x8ec4 */;
                9138: data_o = 32'h00000000 /* 0x8ec8 */;
                9139: data_o = 32'h00000000 /* 0x8ecc */;
                9140: data_o = 32'h00000000 /* 0x8ed0 */;
                9141: data_o = 32'h00000000 /* 0x8ed4 */;
                9142: data_o = 32'h00000000 /* 0x8ed8 */;
                9143: data_o = 32'h00000000 /* 0x8edc */;
                9144: data_o = 32'h00000000 /* 0x8ee0 */;
                9145: data_o = 32'h00000000 /* 0x8ee4 */;
                9146: data_o = 32'h00000000 /* 0x8ee8 */;
                9147: data_o = 32'h00000000 /* 0x8eec */;
                9148: data_o = 32'h00000000 /* 0x8ef0 */;
                9149: data_o = 32'h00000000 /* 0x8ef4 */;
                9150: data_o = 32'h00000000 /* 0x8ef8 */;
                9151: data_o = 32'h00000000 /* 0x8efc */;
                9152: data_o = 32'h00000000 /* 0x8f00 */;
                9153: data_o = 32'h00000000 /* 0x8f04 */;
                9154: data_o = 32'h00000000 /* 0x8f08 */;
                9155: data_o = 32'h00000000 /* 0x8f0c */;
                9156: data_o = 32'h00000000 /* 0x8f10 */;
                9157: data_o = 32'h00000000 /* 0x8f14 */;
                9158: data_o = 32'h00000000 /* 0x8f18 */;
                9159: data_o = 32'h00000000 /* 0x8f1c */;
                9160: data_o = 32'h00000000 /* 0x8f20 */;
                9161: data_o = 32'h00000000 /* 0x8f24 */;
                9162: data_o = 32'h00000000 /* 0x8f28 */;
                9163: data_o = 32'h00000000 /* 0x8f2c */;
                9164: data_o = 32'h00000000 /* 0x8f30 */;
                9165: data_o = 32'h00000000 /* 0x8f34 */;
                9166: data_o = 32'h00000000 /* 0x8f38 */;
                9167: data_o = 32'h00000000 /* 0x8f3c */;
                9168: data_o = 32'h00000000 /* 0x8f40 */;
                9169: data_o = 32'h00000000 /* 0x8f44 */;
                9170: data_o = 32'h00000000 /* 0x8f48 */;
                9171: data_o = 32'h00000000 /* 0x8f4c */;
                9172: data_o = 32'h00000000 /* 0x8f50 */;
                9173: data_o = 32'h00000000 /* 0x8f54 */;
                9174: data_o = 32'h00000000 /* 0x8f58 */;
                9175: data_o = 32'h00000000 /* 0x8f5c */;
                9176: data_o = 32'h00000000 /* 0x8f60 */;
                9177: data_o = 32'h00000000 /* 0x8f64 */;
                9178: data_o = 32'h00000000 /* 0x8f68 */;
                9179: data_o = 32'h00000000 /* 0x8f6c */;
                9180: data_o = 32'h00000000 /* 0x8f70 */;
                9181: data_o = 32'h00000000 /* 0x8f74 */;
                9182: data_o = 32'h00000000 /* 0x8f78 */;
                9183: data_o = 32'h00000000 /* 0x8f7c */;
                9184: data_o = 32'h00000000 /* 0x8f80 */;
                9185: data_o = 32'h00000000 /* 0x8f84 */;
                9186: data_o = 32'h00000000 /* 0x8f88 */;
                9187: data_o = 32'h00000000 /* 0x8f8c */;
                9188: data_o = 32'h00000000 /* 0x8f90 */;
                9189: data_o = 32'h00000000 /* 0x8f94 */;
                9190: data_o = 32'h00000000 /* 0x8f98 */;
                9191: data_o = 32'h00000000 /* 0x8f9c */;
                9192: data_o = 32'h00000000 /* 0x8fa0 */;
                9193: data_o = 32'h00000000 /* 0x8fa4 */;
                9194: data_o = 32'h00000000 /* 0x8fa8 */;
                9195: data_o = 32'h00000000 /* 0x8fac */;
                9196: data_o = 32'h00000000 /* 0x8fb0 */;
                9197: data_o = 32'h00000000 /* 0x8fb4 */;
                9198: data_o = 32'h00000000 /* 0x8fb8 */;
                9199: data_o = 32'h00000000 /* 0x8fbc */;
                9200: data_o = 32'h00000000 /* 0x8fc0 */;
                9201: data_o = 32'h00000000 /* 0x8fc4 */;
                9202: data_o = 32'h00000000 /* 0x8fc8 */;
                9203: data_o = 32'h00000000 /* 0x8fcc */;
                9204: data_o = 32'h00000000 /* 0x8fd0 */;
                9205: data_o = 32'h00000000 /* 0x8fd4 */;
                9206: data_o = 32'h00000000 /* 0x8fd8 */;
                9207: data_o = 32'h00000000 /* 0x8fdc */;
                9208: data_o = 32'h00000000 /* 0x8fe0 */;
                9209: data_o = 32'h00000000 /* 0x8fe4 */;
                9210: data_o = 32'h00000000 /* 0x8fe8 */;
                9211: data_o = 32'h00000000 /* 0x8fec */;
                9212: data_o = 32'h00000000 /* 0x8ff0 */;
                9213: data_o = 32'h00000000 /* 0x8ff4 */;
                9214: data_o = 32'h00000000 /* 0x8ff8 */;
                9215: data_o = 32'h00000000 /* 0x8ffc */;
                9216: data_o = 32'h00000000 /* 0x9000 */;
                9217: data_o = 32'h00000000 /* 0x9004 */;
                9218: data_o = 32'h00000000 /* 0x9008 */;
                9219: data_o = 32'h00000000 /* 0x900c */;
                9220: data_o = 32'h00000000 /* 0x9010 */;
                9221: data_o = 32'h00000000 /* 0x9014 */;
                9222: data_o = 32'h00000000 /* 0x9018 */;
                9223: data_o = 32'h00000000 /* 0x901c */;
                9224: data_o = 32'h00000000 /* 0x9020 */;
                9225: data_o = 32'h00000000 /* 0x9024 */;
                9226: data_o = 32'h00000000 /* 0x9028 */;
                9227: data_o = 32'h00000000 /* 0x902c */;
                9228: data_o = 32'h00000000 /* 0x9030 */;
                9229: data_o = 32'h00000000 /* 0x9034 */;
                9230: data_o = 32'h00000000 /* 0x9038 */;
                9231: data_o = 32'h00000000 /* 0x903c */;
                9232: data_o = 32'h00000000 /* 0x9040 */;
                9233: data_o = 32'h00000000 /* 0x9044 */;
                9234: data_o = 32'h00000000 /* 0x9048 */;
                9235: data_o = 32'h00000000 /* 0x904c */;
                9236: data_o = 32'h00000000 /* 0x9050 */;
                9237: data_o = 32'h00000000 /* 0x9054 */;
                9238: data_o = 32'h00000000 /* 0x9058 */;
                9239: data_o = 32'h00000000 /* 0x905c */;
                9240: data_o = 32'h00000000 /* 0x9060 */;
                9241: data_o = 32'h00000000 /* 0x9064 */;
                9242: data_o = 32'h00000000 /* 0x9068 */;
                9243: data_o = 32'h00000000 /* 0x906c */;
                9244: data_o = 32'h00000000 /* 0x9070 */;
                9245: data_o = 32'h00000000 /* 0x9074 */;
                9246: data_o = 32'h00000000 /* 0x9078 */;
                9247: data_o = 32'h00000000 /* 0x907c */;
                9248: data_o = 32'h00000000 /* 0x9080 */;
                9249: data_o = 32'h00000000 /* 0x9084 */;
                9250: data_o = 32'h00000000 /* 0x9088 */;
                9251: data_o = 32'h00000000 /* 0x908c */;
                9252: data_o = 32'h00000000 /* 0x9090 */;
                9253: data_o = 32'h00000000 /* 0x9094 */;
                9254: data_o = 32'h00000000 /* 0x9098 */;
                9255: data_o = 32'h00000000 /* 0x909c */;
                9256: data_o = 32'h00000000 /* 0x90a0 */;
                9257: data_o = 32'h00000000 /* 0x90a4 */;
                9258: data_o = 32'h00000000 /* 0x90a8 */;
                9259: data_o = 32'h00000000 /* 0x90ac */;
                9260: data_o = 32'h00000000 /* 0x90b0 */;
                9261: data_o = 32'h00000000 /* 0x90b4 */;
                9262: data_o = 32'h00000000 /* 0x90b8 */;
                9263: data_o = 32'h00000000 /* 0x90bc */;
                9264: data_o = 32'h00000000 /* 0x90c0 */;
                9265: data_o = 32'h00000000 /* 0x90c4 */;
                9266: data_o = 32'h00000000 /* 0x90c8 */;
                9267: data_o = 32'h00000000 /* 0x90cc */;
                9268: data_o = 32'h00000000 /* 0x90d0 */;
                9269: data_o = 32'h00000000 /* 0x90d4 */;
                9270: data_o = 32'h00000000 /* 0x90d8 */;
                9271: data_o = 32'h00000000 /* 0x90dc */;
                9272: data_o = 32'h00000000 /* 0x90e0 */;
                9273: data_o = 32'h00000000 /* 0x90e4 */;
                9274: data_o = 32'h00000000 /* 0x90e8 */;
                9275: data_o = 32'h00000000 /* 0x90ec */;
                9276: data_o = 32'h00000000 /* 0x90f0 */;
                9277: data_o = 32'h00000000 /* 0x90f4 */;
                9278: data_o = 32'h00000000 /* 0x90f8 */;
                9279: data_o = 32'h00000000 /* 0x90fc */;
                9280: data_o = 32'h00000000 /* 0x9100 */;
                9281: data_o = 32'h00000000 /* 0x9104 */;
                9282: data_o = 32'h00000000 /* 0x9108 */;
                9283: data_o = 32'h00000000 /* 0x910c */;
                9284: data_o = 32'h00000000 /* 0x9110 */;
                9285: data_o = 32'h00000000 /* 0x9114 */;
                9286: data_o = 32'h00000000 /* 0x9118 */;
                9287: data_o = 32'h00000000 /* 0x911c */;
                9288: data_o = 32'h00000000 /* 0x9120 */;
                9289: data_o = 32'h00000000 /* 0x9124 */;
                9290: data_o = 32'h00000000 /* 0x9128 */;
                9291: data_o = 32'h00000000 /* 0x912c */;
                9292: data_o = 32'h00000000 /* 0x9130 */;
                9293: data_o = 32'h00000000 /* 0x9134 */;
                9294: data_o = 32'h00000000 /* 0x9138 */;
                9295: data_o = 32'h00000000 /* 0x913c */;
                9296: data_o = 32'h00000000 /* 0x9140 */;
                9297: data_o = 32'h00000000 /* 0x9144 */;
                9298: data_o = 32'h00000000 /* 0x9148 */;
                9299: data_o = 32'h00000000 /* 0x914c */;
                9300: data_o = 32'h00000000 /* 0x9150 */;
                9301: data_o = 32'h00000000 /* 0x9154 */;
                9302: data_o = 32'h00000000 /* 0x9158 */;
                9303: data_o = 32'h00000000 /* 0x915c */;
                9304: data_o = 32'h00000000 /* 0x9160 */;
                9305: data_o = 32'h00000000 /* 0x9164 */;
                9306: data_o = 32'h00000000 /* 0x9168 */;
                9307: data_o = 32'h00000000 /* 0x916c */;
                9308: data_o = 32'h00000000 /* 0x9170 */;
                9309: data_o = 32'h00000000 /* 0x9174 */;
                9310: data_o = 32'h00000000 /* 0x9178 */;
                9311: data_o = 32'h00000000 /* 0x917c */;
                9312: data_o = 32'h00000000 /* 0x9180 */;
                9313: data_o = 32'h00000000 /* 0x9184 */;
                9314: data_o = 32'h00000000 /* 0x9188 */;
                9315: data_o = 32'h00000000 /* 0x918c */;
                9316: data_o = 32'h00000000 /* 0x9190 */;
                9317: data_o = 32'h00000000 /* 0x9194 */;
                9318: data_o = 32'h00000000 /* 0x9198 */;
                9319: data_o = 32'h00000000 /* 0x919c */;
                9320: data_o = 32'h00000000 /* 0x91a0 */;
                9321: data_o = 32'h00000000 /* 0x91a4 */;
                9322: data_o = 32'h00000000 /* 0x91a8 */;
                9323: data_o = 32'h00000000 /* 0x91ac */;
                9324: data_o = 32'h00000000 /* 0x91b0 */;
                9325: data_o = 32'h00000000 /* 0x91b4 */;
                9326: data_o = 32'h00000000 /* 0x91b8 */;
                9327: data_o = 32'h00000000 /* 0x91bc */;
                9328: data_o = 32'h00000000 /* 0x91c0 */;
                9329: data_o = 32'h00000000 /* 0x91c4 */;
                9330: data_o = 32'h00000000 /* 0x91c8 */;
                9331: data_o = 32'h00000000 /* 0x91cc */;
                9332: data_o = 32'h00000000 /* 0x91d0 */;
                9333: data_o = 32'h00000000 /* 0x91d4 */;
                9334: data_o = 32'h00000000 /* 0x91d8 */;
                9335: data_o = 32'h00000000 /* 0x91dc */;
                9336: data_o = 32'h00000000 /* 0x91e0 */;
                9337: data_o = 32'h00000000 /* 0x91e4 */;
                9338: data_o = 32'h00000000 /* 0x91e8 */;
                9339: data_o = 32'h00000000 /* 0x91ec */;
                9340: data_o = 32'h00000000 /* 0x91f0 */;
                9341: data_o = 32'h00000000 /* 0x91f4 */;
                9342: data_o = 32'h00000000 /* 0x91f8 */;
                9343: data_o = 32'h00000000 /* 0x91fc */;
                9344: data_o = 32'h00000000 /* 0x9200 */;
                9345: data_o = 32'h00000000 /* 0x9204 */;
                9346: data_o = 32'h00000000 /* 0x9208 */;
                9347: data_o = 32'h00000000 /* 0x920c */;
                9348: data_o = 32'h00000000 /* 0x9210 */;
                9349: data_o = 32'h00000000 /* 0x9214 */;
                9350: data_o = 32'h00000000 /* 0x9218 */;
                9351: data_o = 32'h00000000 /* 0x921c */;
                9352: data_o = 32'h00000000 /* 0x9220 */;
                9353: data_o = 32'h00000000 /* 0x9224 */;
                9354: data_o = 32'h00000000 /* 0x9228 */;
                9355: data_o = 32'h00000000 /* 0x922c */;
                9356: data_o = 32'h00000000 /* 0x9230 */;
                9357: data_o = 32'h00000000 /* 0x9234 */;
                9358: data_o = 32'h00000000 /* 0x9238 */;
                9359: data_o = 32'h00000000 /* 0x923c */;
                9360: data_o = 32'h00000000 /* 0x9240 */;
                9361: data_o = 32'h00000000 /* 0x9244 */;
                9362: data_o = 32'h00000000 /* 0x9248 */;
                9363: data_o = 32'h00000000 /* 0x924c */;
                9364: data_o = 32'h00000000 /* 0x9250 */;
                9365: data_o = 32'h00000000 /* 0x9254 */;
                9366: data_o = 32'h00000000 /* 0x9258 */;
                9367: data_o = 32'h00000000 /* 0x925c */;
                9368: data_o = 32'h00000000 /* 0x9260 */;
                9369: data_o = 32'h00000000 /* 0x9264 */;
                9370: data_o = 32'h00000000 /* 0x9268 */;
                9371: data_o = 32'h00000000 /* 0x926c */;
                9372: data_o = 32'h00000000 /* 0x9270 */;
                9373: data_o = 32'h00000000 /* 0x9274 */;
                9374: data_o = 32'h00000000 /* 0x9278 */;
                9375: data_o = 32'h00000000 /* 0x927c */;
                9376: data_o = 32'h00000000 /* 0x9280 */;
                9377: data_o = 32'h00000000 /* 0x9284 */;
                9378: data_o = 32'h00000000 /* 0x9288 */;
                9379: data_o = 32'h00000000 /* 0x928c */;
                9380: data_o = 32'h00000000 /* 0x9290 */;
                9381: data_o = 32'h00000000 /* 0x9294 */;
                9382: data_o = 32'h00000000 /* 0x9298 */;
                9383: data_o = 32'h00000000 /* 0x929c */;
                9384: data_o = 32'h00000000 /* 0x92a0 */;
                9385: data_o = 32'h00000000 /* 0x92a4 */;
                9386: data_o = 32'h00000000 /* 0x92a8 */;
                9387: data_o = 32'h00000000 /* 0x92ac */;
                9388: data_o = 32'h00000000 /* 0x92b0 */;
                9389: data_o = 32'h00000000 /* 0x92b4 */;
                9390: data_o = 32'h00000000 /* 0x92b8 */;
                9391: data_o = 32'h00000000 /* 0x92bc */;
                9392: data_o = 32'h00000000 /* 0x92c0 */;
                9393: data_o = 32'h00000000 /* 0x92c4 */;
                9394: data_o = 32'h00000000 /* 0x92c8 */;
                9395: data_o = 32'h00000000 /* 0x92cc */;
                9396: data_o = 32'h00000000 /* 0x92d0 */;
                9397: data_o = 32'h00000000 /* 0x92d4 */;
                9398: data_o = 32'h00000000 /* 0x92d8 */;
                9399: data_o = 32'h00000000 /* 0x92dc */;
                9400: data_o = 32'h00000000 /* 0x92e0 */;
                9401: data_o = 32'h00000000 /* 0x92e4 */;
                9402: data_o = 32'h00000000 /* 0x92e8 */;
                9403: data_o = 32'h00000000 /* 0x92ec */;
                9404: data_o = 32'h00000000 /* 0x92f0 */;
                9405: data_o = 32'h00000000 /* 0x92f4 */;
                9406: data_o = 32'h00000000 /* 0x92f8 */;
                9407: data_o = 32'h00000000 /* 0x92fc */;
                9408: data_o = 32'h00000000 /* 0x9300 */;
                9409: data_o = 32'h00000000 /* 0x9304 */;
                9410: data_o = 32'h00000000 /* 0x9308 */;
                9411: data_o = 32'h00000000 /* 0x930c */;
                9412: data_o = 32'h00000000 /* 0x9310 */;
                9413: data_o = 32'h00000000 /* 0x9314 */;
                9414: data_o = 32'h00000000 /* 0x9318 */;
                9415: data_o = 32'h00000000 /* 0x931c */;
                9416: data_o = 32'h00000000 /* 0x9320 */;
                9417: data_o = 32'h00000000 /* 0x9324 */;
                9418: data_o = 32'h00000000 /* 0x9328 */;
                9419: data_o = 32'h00000000 /* 0x932c */;
                9420: data_o = 32'h00000000 /* 0x9330 */;
                9421: data_o = 32'h00000000 /* 0x9334 */;
                9422: data_o = 32'h00000000 /* 0x9338 */;
                9423: data_o = 32'h00000000 /* 0x933c */;
                9424: data_o = 32'h00000000 /* 0x9340 */;
                9425: data_o = 32'h00000000 /* 0x9344 */;
                9426: data_o = 32'h00000000 /* 0x9348 */;
                9427: data_o = 32'h00000000 /* 0x934c */;
                9428: data_o = 32'h00000000 /* 0x9350 */;
                9429: data_o = 32'h00000000 /* 0x9354 */;
                9430: data_o = 32'h00000000 /* 0x9358 */;
                9431: data_o = 32'h00000000 /* 0x935c */;
                9432: data_o = 32'h00000000 /* 0x9360 */;
                9433: data_o = 32'h00000000 /* 0x9364 */;
                9434: data_o = 32'h00000000 /* 0x9368 */;
                9435: data_o = 32'h00000000 /* 0x936c */;
                9436: data_o = 32'h00000000 /* 0x9370 */;
                9437: data_o = 32'h00000000 /* 0x9374 */;
                9438: data_o = 32'h00000000 /* 0x9378 */;
                9439: data_o = 32'h00000000 /* 0x937c */;
                9440: data_o = 32'h00000000 /* 0x9380 */;
                9441: data_o = 32'h00000000 /* 0x9384 */;
                9442: data_o = 32'h00000000 /* 0x9388 */;
                9443: data_o = 32'h00000000 /* 0x938c */;
                9444: data_o = 32'h00000000 /* 0x9390 */;
                9445: data_o = 32'h00000000 /* 0x9394 */;
                9446: data_o = 32'h00000000 /* 0x9398 */;
                9447: data_o = 32'h00000000 /* 0x939c */;
                9448: data_o = 32'h00000000 /* 0x93a0 */;
                9449: data_o = 32'h00000000 /* 0x93a4 */;
                9450: data_o = 32'h00000000 /* 0x93a8 */;
                9451: data_o = 32'h00000000 /* 0x93ac */;
                9452: data_o = 32'h00000000 /* 0x93b0 */;
                9453: data_o = 32'h00000000 /* 0x93b4 */;
                9454: data_o = 32'h00000000 /* 0x93b8 */;
                9455: data_o = 32'h00000000 /* 0x93bc */;
                9456: data_o = 32'h00000000 /* 0x93c0 */;
                9457: data_o = 32'h00000000 /* 0x93c4 */;
                9458: data_o = 32'h00000000 /* 0x93c8 */;
                9459: data_o = 32'h00000000 /* 0x93cc */;
                9460: data_o = 32'h00000000 /* 0x93d0 */;
                9461: data_o = 32'h00000000 /* 0x93d4 */;
                9462: data_o = 32'h00000000 /* 0x93d8 */;
                9463: data_o = 32'h00000000 /* 0x93dc */;
                9464: data_o = 32'h00000000 /* 0x93e0 */;
                9465: data_o = 32'h00000000 /* 0x93e4 */;
                9466: data_o = 32'h00000000 /* 0x93e8 */;
                9467: data_o = 32'h00000000 /* 0x93ec */;
                9468: data_o = 32'h00000000 /* 0x93f0 */;
                9469: data_o = 32'h00000000 /* 0x93f4 */;
                9470: data_o = 32'h00000000 /* 0x93f8 */;
                9471: data_o = 32'h00000000 /* 0x93fc */;
                9472: data_o = 32'h00000000 /* 0x9400 */;
                9473: data_o = 32'h00000000 /* 0x9404 */;
                9474: data_o = 32'h00000000 /* 0x9408 */;
                9475: data_o = 32'h00000000 /* 0x940c */;
                9476: data_o = 32'h00000000 /* 0x9410 */;
                9477: data_o = 32'h00000000 /* 0x9414 */;
                9478: data_o = 32'h00000000 /* 0x9418 */;
                9479: data_o = 32'h00000000 /* 0x941c */;
                9480: data_o = 32'h00000000 /* 0x9420 */;
                9481: data_o = 32'h00000000 /* 0x9424 */;
                9482: data_o = 32'h00000000 /* 0x9428 */;
                9483: data_o = 32'h00000000 /* 0x942c */;
                9484: data_o = 32'h00000000 /* 0x9430 */;
                9485: data_o = 32'h00000000 /* 0x9434 */;
                9486: data_o = 32'h00000000 /* 0x9438 */;
                9487: data_o = 32'h00000000 /* 0x943c */;
                9488: data_o = 32'h00000000 /* 0x9440 */;
                9489: data_o = 32'h00000000 /* 0x9444 */;
                9490: data_o = 32'h00000000 /* 0x9448 */;
                9491: data_o = 32'h00000000 /* 0x944c */;
                9492: data_o = 32'h00000000 /* 0x9450 */;
                9493: data_o = 32'h00000000 /* 0x9454 */;
                9494: data_o = 32'h00000000 /* 0x9458 */;
                9495: data_o = 32'h00000000 /* 0x945c */;
                9496: data_o = 32'h00000000 /* 0x9460 */;
                9497: data_o = 32'h00000000 /* 0x9464 */;
                9498: data_o = 32'h00000000 /* 0x9468 */;
                9499: data_o = 32'h00000000 /* 0x946c */;
                9500: data_o = 32'h00000000 /* 0x9470 */;
                9501: data_o = 32'h00000000 /* 0x9474 */;
                9502: data_o = 32'h00000000 /* 0x9478 */;
                9503: data_o = 32'h00000000 /* 0x947c */;
                9504: data_o = 32'h00000000 /* 0x9480 */;
                9505: data_o = 32'h00000000 /* 0x9484 */;
                9506: data_o = 32'h00000000 /* 0x9488 */;
                9507: data_o = 32'h00000000 /* 0x948c */;
                9508: data_o = 32'h00000000 /* 0x9490 */;
                9509: data_o = 32'h00000000 /* 0x9494 */;
                9510: data_o = 32'h00000000 /* 0x9498 */;
                9511: data_o = 32'h00000000 /* 0x949c */;
                9512: data_o = 32'h00000000 /* 0x94a0 */;
                9513: data_o = 32'h00000000 /* 0x94a4 */;
                9514: data_o = 32'h00000000 /* 0x94a8 */;
                9515: data_o = 32'h00000000 /* 0x94ac */;
                9516: data_o = 32'h00000000 /* 0x94b0 */;
                9517: data_o = 32'h00000000 /* 0x94b4 */;
                9518: data_o = 32'h00000000 /* 0x94b8 */;
                9519: data_o = 32'h00000000 /* 0x94bc */;
                9520: data_o = 32'h00000000 /* 0x94c0 */;
                9521: data_o = 32'h00000000 /* 0x94c4 */;
                9522: data_o = 32'h00000000 /* 0x94c8 */;
                9523: data_o = 32'h00000000 /* 0x94cc */;
                9524: data_o = 32'h00000000 /* 0x94d0 */;
                9525: data_o = 32'h00000000 /* 0x94d4 */;
                9526: data_o = 32'h00000000 /* 0x94d8 */;
                9527: data_o = 32'h00000000 /* 0x94dc */;
                9528: data_o = 32'h00000000 /* 0x94e0 */;
                9529: data_o = 32'h00000000 /* 0x94e4 */;
                9530: data_o = 32'h00000000 /* 0x94e8 */;
                9531: data_o = 32'h00000000 /* 0x94ec */;
                9532: data_o = 32'h00000000 /* 0x94f0 */;
                9533: data_o = 32'h00000000 /* 0x94f4 */;
                9534: data_o = 32'h00000000 /* 0x94f8 */;
                9535: data_o = 32'h00000000 /* 0x94fc */;
                9536: data_o = 32'h00000000 /* 0x9500 */;
                9537: data_o = 32'h00000000 /* 0x9504 */;
                9538: data_o = 32'h00000000 /* 0x9508 */;
                9539: data_o = 32'h00000000 /* 0x950c */;
                9540: data_o = 32'h00000000 /* 0x9510 */;
                9541: data_o = 32'h00000000 /* 0x9514 */;
                9542: data_o = 32'h00000000 /* 0x9518 */;
                9543: data_o = 32'h00000000 /* 0x951c */;
                9544: data_o = 32'h00000000 /* 0x9520 */;
                9545: data_o = 32'h00000000 /* 0x9524 */;
                9546: data_o = 32'h00000000 /* 0x9528 */;
                9547: data_o = 32'h00000000 /* 0x952c */;
                9548: data_o = 32'h00000000 /* 0x9530 */;
                9549: data_o = 32'h00000000 /* 0x9534 */;
                9550: data_o = 32'h00000000 /* 0x9538 */;
                9551: data_o = 32'h00000000 /* 0x953c */;
                9552: data_o = 32'h00000000 /* 0x9540 */;
                9553: data_o = 32'h00000000 /* 0x9544 */;
                9554: data_o = 32'h00000000 /* 0x9548 */;
                9555: data_o = 32'h00000000 /* 0x954c */;
                9556: data_o = 32'h00000000 /* 0x9550 */;
                9557: data_o = 32'h00000000 /* 0x9554 */;
                9558: data_o = 32'h00000000 /* 0x9558 */;
                9559: data_o = 32'h00000000 /* 0x955c */;
                9560: data_o = 32'h00000000 /* 0x9560 */;
                9561: data_o = 32'h00000000 /* 0x9564 */;
                9562: data_o = 32'h00000000 /* 0x9568 */;
                9563: data_o = 32'h00000000 /* 0x956c */;
                9564: data_o = 32'h00000000 /* 0x9570 */;
                9565: data_o = 32'h00000000 /* 0x9574 */;
                9566: data_o = 32'h00000000 /* 0x9578 */;
                9567: data_o = 32'h00000000 /* 0x957c */;
                9568: data_o = 32'h00000000 /* 0x9580 */;
                9569: data_o = 32'h00000000 /* 0x9584 */;
                9570: data_o = 32'h00000000 /* 0x9588 */;
                9571: data_o = 32'h00000000 /* 0x958c */;
                9572: data_o = 32'h00000000 /* 0x9590 */;
                9573: data_o = 32'h00000000 /* 0x9594 */;
                9574: data_o = 32'h00000000 /* 0x9598 */;
                9575: data_o = 32'h00000000 /* 0x959c */;
                9576: data_o = 32'h00000000 /* 0x95a0 */;
                9577: data_o = 32'h00000000 /* 0x95a4 */;
                9578: data_o = 32'h00000000 /* 0x95a8 */;
                9579: data_o = 32'h00000000 /* 0x95ac */;
                9580: data_o = 32'h00000000 /* 0x95b0 */;
                9581: data_o = 32'h00000000 /* 0x95b4 */;
                9582: data_o = 32'h00000000 /* 0x95b8 */;
                9583: data_o = 32'h00000000 /* 0x95bc */;
                9584: data_o = 32'h00000000 /* 0x95c0 */;
                9585: data_o = 32'h00000000 /* 0x95c4 */;
                9586: data_o = 32'h00000000 /* 0x95c8 */;
                9587: data_o = 32'h00000000 /* 0x95cc */;
                9588: data_o = 32'h00000000 /* 0x95d0 */;
                9589: data_o = 32'h00000000 /* 0x95d4 */;
                9590: data_o = 32'h00000000 /* 0x95d8 */;
                9591: data_o = 32'h00000000 /* 0x95dc */;
                9592: data_o = 32'h00000000 /* 0x95e0 */;
                9593: data_o = 32'h00000000 /* 0x95e4 */;
                9594: data_o = 32'h00000000 /* 0x95e8 */;
                9595: data_o = 32'h00000000 /* 0x95ec */;
                9596: data_o = 32'h00000000 /* 0x95f0 */;
                9597: data_o = 32'h00000000 /* 0x95f4 */;
                9598: data_o = 32'h00000000 /* 0x95f8 */;
                9599: data_o = 32'h00000000 /* 0x95fc */;
                9600: data_o = 32'h00000000 /* 0x9600 */;
                9601: data_o = 32'h00000000 /* 0x9604 */;
                9602: data_o = 32'h00000000 /* 0x9608 */;
                9603: data_o = 32'h00000000 /* 0x960c */;
                9604: data_o = 32'h00000000 /* 0x9610 */;
                9605: data_o = 32'h00000000 /* 0x9614 */;
                9606: data_o = 32'h00000000 /* 0x9618 */;
                9607: data_o = 32'h00000000 /* 0x961c */;
                9608: data_o = 32'h00000000 /* 0x9620 */;
                9609: data_o = 32'h00000000 /* 0x9624 */;
                9610: data_o = 32'h00000000 /* 0x9628 */;
                9611: data_o = 32'h00000000 /* 0x962c */;
                9612: data_o = 32'h00000000 /* 0x9630 */;
                9613: data_o = 32'h00000000 /* 0x9634 */;
                9614: data_o = 32'h00000000 /* 0x9638 */;
                9615: data_o = 32'h00000000 /* 0x963c */;
                9616: data_o = 32'h00000000 /* 0x9640 */;
                9617: data_o = 32'h00000000 /* 0x9644 */;
                9618: data_o = 32'h00000000 /* 0x9648 */;
                9619: data_o = 32'h00000000 /* 0x964c */;
                9620: data_o = 32'h00000000 /* 0x9650 */;
                9621: data_o = 32'h00000000 /* 0x9654 */;
                9622: data_o = 32'h00000000 /* 0x9658 */;
                9623: data_o = 32'h00000000 /* 0x965c */;
                9624: data_o = 32'h00000000 /* 0x9660 */;
                9625: data_o = 32'h00000000 /* 0x9664 */;
                9626: data_o = 32'h00000000 /* 0x9668 */;
                9627: data_o = 32'h00000000 /* 0x966c */;
                9628: data_o = 32'h00000000 /* 0x9670 */;
                9629: data_o = 32'h00000000 /* 0x9674 */;
                9630: data_o = 32'h00000000 /* 0x9678 */;
                9631: data_o = 32'h00000000 /* 0x967c */;
                9632: data_o = 32'h00000000 /* 0x9680 */;
                9633: data_o = 32'h00000000 /* 0x9684 */;
                9634: data_o = 32'h00000000 /* 0x9688 */;
                9635: data_o = 32'h00000000 /* 0x968c */;
                9636: data_o = 32'h00000000 /* 0x9690 */;
                9637: data_o = 32'h00000000 /* 0x9694 */;
                9638: data_o = 32'h00000000 /* 0x9698 */;
                9639: data_o = 32'h00000000 /* 0x969c */;
                9640: data_o = 32'h00000000 /* 0x96a0 */;
                9641: data_o = 32'h00000000 /* 0x96a4 */;
                9642: data_o = 32'h00000000 /* 0x96a8 */;
                9643: data_o = 32'h00000000 /* 0x96ac */;
                9644: data_o = 32'h00000000 /* 0x96b0 */;
                9645: data_o = 32'h00000000 /* 0x96b4 */;
                9646: data_o = 32'h00000000 /* 0x96b8 */;
                9647: data_o = 32'h00000000 /* 0x96bc */;
                9648: data_o = 32'h00000000 /* 0x96c0 */;
                9649: data_o = 32'h00000000 /* 0x96c4 */;
                9650: data_o = 32'h00000000 /* 0x96c8 */;
                9651: data_o = 32'h00000000 /* 0x96cc */;
                9652: data_o = 32'h00000000 /* 0x96d0 */;
                9653: data_o = 32'h00000000 /* 0x96d4 */;
                9654: data_o = 32'h00000000 /* 0x96d8 */;
                9655: data_o = 32'h00000000 /* 0x96dc */;
                9656: data_o = 32'h00000000 /* 0x96e0 */;
                9657: data_o = 32'h00000000 /* 0x96e4 */;
                9658: data_o = 32'h00000000 /* 0x96e8 */;
                9659: data_o = 32'h00000000 /* 0x96ec */;
                9660: data_o = 32'h00000000 /* 0x96f0 */;
                9661: data_o = 32'h00000000 /* 0x96f4 */;
                9662: data_o = 32'h00000000 /* 0x96f8 */;
                9663: data_o = 32'h00000000 /* 0x96fc */;
                9664: data_o = 32'h00000000 /* 0x9700 */;
                9665: data_o = 32'h00000000 /* 0x9704 */;
                9666: data_o = 32'h00000000 /* 0x9708 */;
                9667: data_o = 32'h00000000 /* 0x970c */;
                9668: data_o = 32'h00000000 /* 0x9710 */;
                9669: data_o = 32'h00000000 /* 0x9714 */;
                9670: data_o = 32'h00000000 /* 0x9718 */;
                9671: data_o = 32'h00000000 /* 0x971c */;
                9672: data_o = 32'h00000000 /* 0x9720 */;
                9673: data_o = 32'h00000000 /* 0x9724 */;
                9674: data_o = 32'h00000000 /* 0x9728 */;
                9675: data_o = 32'h00000000 /* 0x972c */;
                9676: data_o = 32'h00000000 /* 0x9730 */;
                9677: data_o = 32'h00000000 /* 0x9734 */;
                9678: data_o = 32'h00000000 /* 0x9738 */;
                9679: data_o = 32'h00000000 /* 0x973c */;
                9680: data_o = 32'h00000000 /* 0x9740 */;
                9681: data_o = 32'h00000000 /* 0x9744 */;
                9682: data_o = 32'h00000000 /* 0x9748 */;
                9683: data_o = 32'h00000000 /* 0x974c */;
                9684: data_o = 32'h00000000 /* 0x9750 */;
                9685: data_o = 32'h00000000 /* 0x9754 */;
                9686: data_o = 32'h00000000 /* 0x9758 */;
                9687: data_o = 32'h00000000 /* 0x975c */;
                9688: data_o = 32'h00000000 /* 0x9760 */;
                9689: data_o = 32'h00000000 /* 0x9764 */;
                9690: data_o = 32'h00000000 /* 0x9768 */;
                9691: data_o = 32'h00000000 /* 0x976c */;
                9692: data_o = 32'h00000000 /* 0x9770 */;
                9693: data_o = 32'h00000000 /* 0x9774 */;
                9694: data_o = 32'h00000000 /* 0x9778 */;
                9695: data_o = 32'h00000000 /* 0x977c */;
                9696: data_o = 32'h00000000 /* 0x9780 */;
                9697: data_o = 32'h00000000 /* 0x9784 */;
                9698: data_o = 32'h00000000 /* 0x9788 */;
                9699: data_o = 32'h00000000 /* 0x978c */;
                9700: data_o = 32'h00000000 /* 0x9790 */;
                9701: data_o = 32'h00000000 /* 0x9794 */;
                9702: data_o = 32'h00000000 /* 0x9798 */;
                9703: data_o = 32'h00000000 /* 0x979c */;
                9704: data_o = 32'h00000000 /* 0x97a0 */;
                9705: data_o = 32'h00000000 /* 0x97a4 */;
                9706: data_o = 32'h00000000 /* 0x97a8 */;
                9707: data_o = 32'h00000000 /* 0x97ac */;
                9708: data_o = 32'h00000000 /* 0x97b0 */;
                9709: data_o = 32'h00000000 /* 0x97b4 */;
                9710: data_o = 32'h00000000 /* 0x97b8 */;
                9711: data_o = 32'h00000000 /* 0x97bc */;
                9712: data_o = 32'h00000000 /* 0x97c0 */;
                9713: data_o = 32'h00000000 /* 0x97c4 */;
                9714: data_o = 32'h00000000 /* 0x97c8 */;
                9715: data_o = 32'h00000000 /* 0x97cc */;
                9716: data_o = 32'h00000000 /* 0x97d0 */;
                9717: data_o = 32'h00000000 /* 0x97d4 */;
                9718: data_o = 32'h00000000 /* 0x97d8 */;
                9719: data_o = 32'h00000000 /* 0x97dc */;
                9720: data_o = 32'h00000000 /* 0x97e0 */;
                9721: data_o = 32'h00000000 /* 0x97e4 */;
                9722: data_o = 32'h00000000 /* 0x97e8 */;
                9723: data_o = 32'h00000000 /* 0x97ec */;
                9724: data_o = 32'h00000000 /* 0x97f0 */;
                9725: data_o = 32'h00000000 /* 0x97f4 */;
                9726: data_o = 32'h00000000 /* 0x97f8 */;
                9727: data_o = 32'h00000000 /* 0x97fc */;
                9728: data_o = 32'h00000000 /* 0x9800 */;
                9729: data_o = 32'h00000000 /* 0x9804 */;
                9730: data_o = 32'h00000000 /* 0x9808 */;
                9731: data_o = 32'h00000000 /* 0x980c */;
                9732: data_o = 32'h00000000 /* 0x9810 */;
                9733: data_o = 32'h00000000 /* 0x9814 */;
                9734: data_o = 32'h00000000 /* 0x9818 */;
                9735: data_o = 32'h00000000 /* 0x981c */;
                9736: data_o = 32'h00000000 /* 0x9820 */;
                9737: data_o = 32'h00000000 /* 0x9824 */;
                9738: data_o = 32'h00000000 /* 0x9828 */;
                9739: data_o = 32'h00000000 /* 0x982c */;
                9740: data_o = 32'h00000000 /* 0x9830 */;
                9741: data_o = 32'h00000000 /* 0x9834 */;
                9742: data_o = 32'h00000000 /* 0x9838 */;
                9743: data_o = 32'h00000000 /* 0x983c */;
                9744: data_o = 32'h00000000 /* 0x9840 */;
                9745: data_o = 32'h00000000 /* 0x9844 */;
                9746: data_o = 32'h00000000 /* 0x9848 */;
                9747: data_o = 32'h00000000 /* 0x984c */;
                9748: data_o = 32'h00000000 /* 0x9850 */;
                9749: data_o = 32'h00000000 /* 0x9854 */;
                9750: data_o = 32'h00000000 /* 0x9858 */;
                9751: data_o = 32'h00000000 /* 0x985c */;
                9752: data_o = 32'h00000000 /* 0x9860 */;
                9753: data_o = 32'h00000000 /* 0x9864 */;
                9754: data_o = 32'h00000000 /* 0x9868 */;
                9755: data_o = 32'h00000000 /* 0x986c */;
                9756: data_o = 32'h00000000 /* 0x9870 */;
                9757: data_o = 32'h00000000 /* 0x9874 */;
                9758: data_o = 32'h00000000 /* 0x9878 */;
                9759: data_o = 32'h00000000 /* 0x987c */;
                9760: data_o = 32'h00000000 /* 0x9880 */;
                9761: data_o = 32'h00000000 /* 0x9884 */;
                9762: data_o = 32'h00000000 /* 0x9888 */;
                9763: data_o = 32'h00000000 /* 0x988c */;
                9764: data_o = 32'h00000000 /* 0x9890 */;
                9765: data_o = 32'h00000000 /* 0x9894 */;
                9766: data_o = 32'h00000000 /* 0x9898 */;
                9767: data_o = 32'h00000000 /* 0x989c */;
                9768: data_o = 32'h00000000 /* 0x98a0 */;
                9769: data_o = 32'h00000000 /* 0x98a4 */;
                9770: data_o = 32'h00000000 /* 0x98a8 */;
                9771: data_o = 32'h00000000 /* 0x98ac */;
                9772: data_o = 32'h00000000 /* 0x98b0 */;
                9773: data_o = 32'h00000000 /* 0x98b4 */;
                9774: data_o = 32'h00000000 /* 0x98b8 */;
                9775: data_o = 32'h00000000 /* 0x98bc */;
                9776: data_o = 32'h00000000 /* 0x98c0 */;
                9777: data_o = 32'h00000000 /* 0x98c4 */;
                9778: data_o = 32'h00000000 /* 0x98c8 */;
                9779: data_o = 32'h00000000 /* 0x98cc */;
                9780: data_o = 32'h00000000 /* 0x98d0 */;
                9781: data_o = 32'h00000000 /* 0x98d4 */;
                9782: data_o = 32'h00000000 /* 0x98d8 */;
                9783: data_o = 32'h00000000 /* 0x98dc */;
                9784: data_o = 32'h00000000 /* 0x98e0 */;
                9785: data_o = 32'h00000000 /* 0x98e4 */;
                9786: data_o = 32'h00000000 /* 0x98e8 */;
                9787: data_o = 32'h00000000 /* 0x98ec */;
                9788: data_o = 32'h00000000 /* 0x98f0 */;
                9789: data_o = 32'h00000000 /* 0x98f4 */;
                9790: data_o = 32'h00000000 /* 0x98f8 */;
                9791: data_o = 32'h00000000 /* 0x98fc */;
                9792: data_o = 32'h00000000 /* 0x9900 */;
                9793: data_o = 32'h00000000 /* 0x9904 */;
                9794: data_o = 32'h00000000 /* 0x9908 */;
                9795: data_o = 32'h00000000 /* 0x990c */;
                9796: data_o = 32'h00000000 /* 0x9910 */;
                9797: data_o = 32'h00000000 /* 0x9914 */;
                9798: data_o = 32'h00000000 /* 0x9918 */;
                9799: data_o = 32'h00000000 /* 0x991c */;
                9800: data_o = 32'h00000000 /* 0x9920 */;
                9801: data_o = 32'h00000000 /* 0x9924 */;
                9802: data_o = 32'h00000000 /* 0x9928 */;
                9803: data_o = 32'h00000000 /* 0x992c */;
                9804: data_o = 32'h00000000 /* 0x9930 */;
                9805: data_o = 32'h00000000 /* 0x9934 */;
                9806: data_o = 32'h00000000 /* 0x9938 */;
                9807: data_o = 32'h00000000 /* 0x993c */;
                9808: data_o = 32'h00000000 /* 0x9940 */;
                9809: data_o = 32'h00000000 /* 0x9944 */;
                9810: data_o = 32'h00000000 /* 0x9948 */;
                9811: data_o = 32'h00000000 /* 0x994c */;
                9812: data_o = 32'h00000000 /* 0x9950 */;
                9813: data_o = 32'h00000000 /* 0x9954 */;
                9814: data_o = 32'h00000000 /* 0x9958 */;
                9815: data_o = 32'h00000000 /* 0x995c */;
                9816: data_o = 32'h00000000 /* 0x9960 */;
                9817: data_o = 32'h00000000 /* 0x9964 */;
                9818: data_o = 32'h00000000 /* 0x9968 */;
                9819: data_o = 32'h00000000 /* 0x996c */;
                9820: data_o = 32'h00000000 /* 0x9970 */;
                9821: data_o = 32'h00000000 /* 0x9974 */;
                9822: data_o = 32'h00000000 /* 0x9978 */;
                9823: data_o = 32'h00000000 /* 0x997c */;
                9824: data_o = 32'h00000000 /* 0x9980 */;
                9825: data_o = 32'h00000000 /* 0x9984 */;
                9826: data_o = 32'h00000000 /* 0x9988 */;
                9827: data_o = 32'h00000000 /* 0x998c */;
                9828: data_o = 32'h00000000 /* 0x9990 */;
                9829: data_o = 32'h00000000 /* 0x9994 */;
                9830: data_o = 32'h00000000 /* 0x9998 */;
                9831: data_o = 32'h00000000 /* 0x999c */;
                9832: data_o = 32'h00000000 /* 0x99a0 */;
                9833: data_o = 32'h00000000 /* 0x99a4 */;
                9834: data_o = 32'h00000000 /* 0x99a8 */;
                9835: data_o = 32'h00000000 /* 0x99ac */;
                9836: data_o = 32'h00000000 /* 0x99b0 */;
                9837: data_o = 32'h00000000 /* 0x99b4 */;
                9838: data_o = 32'h00000000 /* 0x99b8 */;
                9839: data_o = 32'h00000000 /* 0x99bc */;
                9840: data_o = 32'h00000000 /* 0x99c0 */;
                9841: data_o = 32'h00000000 /* 0x99c4 */;
                9842: data_o = 32'h00000000 /* 0x99c8 */;
                9843: data_o = 32'h00000000 /* 0x99cc */;
                9844: data_o = 32'h00000000 /* 0x99d0 */;
                9845: data_o = 32'h00000000 /* 0x99d4 */;
                9846: data_o = 32'h00000000 /* 0x99d8 */;
                9847: data_o = 32'h00000000 /* 0x99dc */;
                9848: data_o = 32'h00000000 /* 0x99e0 */;
                9849: data_o = 32'h00000000 /* 0x99e4 */;
                9850: data_o = 32'h00000000 /* 0x99e8 */;
                9851: data_o = 32'h00000000 /* 0x99ec */;
                9852: data_o = 32'h00000000 /* 0x99f0 */;
                9853: data_o = 32'h00000000 /* 0x99f4 */;
                9854: data_o = 32'h00000000 /* 0x99f8 */;
                9855: data_o = 32'h00000000 /* 0x99fc */;
                9856: data_o = 32'h00000000 /* 0x9a00 */;
                9857: data_o = 32'h00000000 /* 0x9a04 */;
                9858: data_o = 32'h00000000 /* 0x9a08 */;
                9859: data_o = 32'h00000000 /* 0x9a0c */;
                9860: data_o = 32'h00000000 /* 0x9a10 */;
                9861: data_o = 32'h00000000 /* 0x9a14 */;
                9862: data_o = 32'h00000000 /* 0x9a18 */;
                9863: data_o = 32'h00000000 /* 0x9a1c */;
                9864: data_o = 32'h00000000 /* 0x9a20 */;
                9865: data_o = 32'h00000000 /* 0x9a24 */;
                9866: data_o = 32'h00000000 /* 0x9a28 */;
                9867: data_o = 32'h00000000 /* 0x9a2c */;
                9868: data_o = 32'h00000000 /* 0x9a30 */;
                9869: data_o = 32'h00000000 /* 0x9a34 */;
                9870: data_o = 32'h00000000 /* 0x9a38 */;
                9871: data_o = 32'h00000000 /* 0x9a3c */;
                9872: data_o = 32'h00000000 /* 0x9a40 */;
                9873: data_o = 32'h00000000 /* 0x9a44 */;
                9874: data_o = 32'h00000000 /* 0x9a48 */;
                9875: data_o = 32'h00000000 /* 0x9a4c */;
                9876: data_o = 32'h00000000 /* 0x9a50 */;
                9877: data_o = 32'h00000000 /* 0x9a54 */;
                9878: data_o = 32'h00000000 /* 0x9a58 */;
                9879: data_o = 32'h00000000 /* 0x9a5c */;
                9880: data_o = 32'h00000000 /* 0x9a60 */;
                9881: data_o = 32'h00000000 /* 0x9a64 */;
                9882: data_o = 32'h00000000 /* 0x9a68 */;
                9883: data_o = 32'h00000000 /* 0x9a6c */;
                9884: data_o = 32'h00000000 /* 0x9a70 */;
                9885: data_o = 32'h00000000 /* 0x9a74 */;
                9886: data_o = 32'h00000000 /* 0x9a78 */;
                9887: data_o = 32'h00000000 /* 0x9a7c */;
                9888: data_o = 32'h00000000 /* 0x9a80 */;
                9889: data_o = 32'h00000000 /* 0x9a84 */;
                9890: data_o = 32'h00000000 /* 0x9a88 */;
                9891: data_o = 32'h00000000 /* 0x9a8c */;
                9892: data_o = 32'h00000000 /* 0x9a90 */;
                9893: data_o = 32'h00000000 /* 0x9a94 */;
                9894: data_o = 32'h00000000 /* 0x9a98 */;
                9895: data_o = 32'h00000000 /* 0x9a9c */;
                9896: data_o = 32'h00000000 /* 0x9aa0 */;
                9897: data_o = 32'h00000000 /* 0x9aa4 */;
                9898: data_o = 32'h00000000 /* 0x9aa8 */;
                9899: data_o = 32'h00000000 /* 0x9aac */;
                9900: data_o = 32'h00000000 /* 0x9ab0 */;
                9901: data_o = 32'h00000000 /* 0x9ab4 */;
                9902: data_o = 32'h00000000 /* 0x9ab8 */;
                9903: data_o = 32'h00000000 /* 0x9abc */;
                9904: data_o = 32'h00000000 /* 0x9ac0 */;
                9905: data_o = 32'h00000000 /* 0x9ac4 */;
                9906: data_o = 32'h00000000 /* 0x9ac8 */;
                9907: data_o = 32'h00000000 /* 0x9acc */;
                9908: data_o = 32'h00000000 /* 0x9ad0 */;
                9909: data_o = 32'h00000000 /* 0x9ad4 */;
                9910: data_o = 32'h00000000 /* 0x9ad8 */;
                9911: data_o = 32'h00000000 /* 0x9adc */;
                9912: data_o = 32'h00000000 /* 0x9ae0 */;
                9913: data_o = 32'h00000000 /* 0x9ae4 */;
                9914: data_o = 32'h00000000 /* 0x9ae8 */;
                9915: data_o = 32'h00000000 /* 0x9aec */;
                9916: data_o = 32'h00000000 /* 0x9af0 */;
                9917: data_o = 32'h00000000 /* 0x9af4 */;
                9918: data_o = 32'h00000000 /* 0x9af8 */;
                9919: data_o = 32'h00000000 /* 0x9afc */;
                9920: data_o = 32'h00000000 /* 0x9b00 */;
                9921: data_o = 32'h00000000 /* 0x9b04 */;
                9922: data_o = 32'h00000000 /* 0x9b08 */;
                9923: data_o = 32'h00000000 /* 0x9b0c */;
                9924: data_o = 32'h00000000 /* 0x9b10 */;
                9925: data_o = 32'h00000000 /* 0x9b14 */;
                9926: data_o = 32'h00000000 /* 0x9b18 */;
                9927: data_o = 32'h00000000 /* 0x9b1c */;
                9928: data_o = 32'h00000000 /* 0x9b20 */;
                9929: data_o = 32'h00000000 /* 0x9b24 */;
                9930: data_o = 32'h00000000 /* 0x9b28 */;
                9931: data_o = 32'h00000000 /* 0x9b2c */;
                9932: data_o = 32'h00000000 /* 0x9b30 */;
                9933: data_o = 32'h00000000 /* 0x9b34 */;
                9934: data_o = 32'h00000000 /* 0x9b38 */;
                9935: data_o = 32'h00000000 /* 0x9b3c */;
                9936: data_o = 32'h00000000 /* 0x9b40 */;
                9937: data_o = 32'h00000000 /* 0x9b44 */;
                9938: data_o = 32'h00000000 /* 0x9b48 */;
                9939: data_o = 32'h00000000 /* 0x9b4c */;
                9940: data_o = 32'h00000000 /* 0x9b50 */;
                9941: data_o = 32'h00000000 /* 0x9b54 */;
                9942: data_o = 32'h00000000 /* 0x9b58 */;
                9943: data_o = 32'h00000000 /* 0x9b5c */;
                9944: data_o = 32'h00000000 /* 0x9b60 */;
                9945: data_o = 32'h00000000 /* 0x9b64 */;
                9946: data_o = 32'h00000000 /* 0x9b68 */;
                9947: data_o = 32'h00000000 /* 0x9b6c */;
                9948: data_o = 32'h00000000 /* 0x9b70 */;
                9949: data_o = 32'h00000000 /* 0x9b74 */;
                9950: data_o = 32'h00000000 /* 0x9b78 */;
                9951: data_o = 32'h00000000 /* 0x9b7c */;
                9952: data_o = 32'h00000000 /* 0x9b80 */;
                9953: data_o = 32'h00000000 /* 0x9b84 */;
                9954: data_o = 32'h00000000 /* 0x9b88 */;
                9955: data_o = 32'h00000000 /* 0x9b8c */;
                9956: data_o = 32'h00000000 /* 0x9b90 */;
                9957: data_o = 32'h00000000 /* 0x9b94 */;
                9958: data_o = 32'h00000000 /* 0x9b98 */;
                9959: data_o = 32'h00000000 /* 0x9b9c */;
                9960: data_o = 32'h00000000 /* 0x9ba0 */;
                9961: data_o = 32'h00000000 /* 0x9ba4 */;
                9962: data_o = 32'h00000000 /* 0x9ba8 */;
                9963: data_o = 32'h00000000 /* 0x9bac */;
                9964: data_o = 32'h00000000 /* 0x9bb0 */;
                9965: data_o = 32'h00000000 /* 0x9bb4 */;
                9966: data_o = 32'h00000000 /* 0x9bb8 */;
                9967: data_o = 32'h00000000 /* 0x9bbc */;
                9968: data_o = 32'h00000000 /* 0x9bc0 */;
                9969: data_o = 32'h00000000 /* 0x9bc4 */;
                9970: data_o = 32'h00000000 /* 0x9bc8 */;
                9971: data_o = 32'h00000000 /* 0x9bcc */;
                9972: data_o = 32'h00000000 /* 0x9bd0 */;
                9973: data_o = 32'h00000000 /* 0x9bd4 */;
                9974: data_o = 32'h00000000 /* 0x9bd8 */;
                9975: data_o = 32'h00000000 /* 0x9bdc */;
                9976: data_o = 32'h00000000 /* 0x9be0 */;
                9977: data_o = 32'h00000000 /* 0x9be4 */;
                9978: data_o = 32'h00000000 /* 0x9be8 */;
                9979: data_o = 32'h00000000 /* 0x9bec */;
                9980: data_o = 32'h00000000 /* 0x9bf0 */;
                9981: data_o = 32'h00000000 /* 0x9bf4 */;
                9982: data_o = 32'h00000000 /* 0x9bf8 */;
                9983: data_o = 32'h00000000 /* 0x9bfc */;
                9984: data_o = 32'h00000000 /* 0x9c00 */;
                9985: data_o = 32'h00000000 /* 0x9c04 */;
                9986: data_o = 32'h00000000 /* 0x9c08 */;
                9987: data_o = 32'h00000000 /* 0x9c0c */;
                9988: data_o = 32'h00000000 /* 0x9c10 */;
                9989: data_o = 32'h00000000 /* 0x9c14 */;
                9990: data_o = 32'h00000000 /* 0x9c18 */;
                9991: data_o = 32'h00000000 /* 0x9c1c */;
                9992: data_o = 32'h00000000 /* 0x9c20 */;
                9993: data_o = 32'h00000000 /* 0x9c24 */;
                9994: data_o = 32'h00000000 /* 0x9c28 */;
                9995: data_o = 32'h00000000 /* 0x9c2c */;
                9996: data_o = 32'h00000000 /* 0x9c30 */;
                9997: data_o = 32'h00000000 /* 0x9c34 */;
                9998: data_o = 32'h00000000 /* 0x9c38 */;
                9999: data_o = 32'h00000000 /* 0x9c3c */;
                10000: data_o = 32'h00000000 /* 0x9c40 */;
                10001: data_o = 32'h00000000 /* 0x9c44 */;
                10002: data_o = 32'h00000000 /* 0x9c48 */;
                10003: data_o = 32'h00000000 /* 0x9c4c */;
                10004: data_o = 32'h00000000 /* 0x9c50 */;
                10005: data_o = 32'h00000000 /* 0x9c54 */;
                10006: data_o = 32'h00000000 /* 0x9c58 */;
                10007: data_o = 32'h00000000 /* 0x9c5c */;
                10008: data_o = 32'h00000000 /* 0x9c60 */;
                10009: data_o = 32'h00000000 /* 0x9c64 */;
                10010: data_o = 32'h00000000 /* 0x9c68 */;
                10011: data_o = 32'h00000000 /* 0x9c6c */;
                10012: data_o = 32'h00000000 /* 0x9c70 */;
                10013: data_o = 32'h00000000 /* 0x9c74 */;
                10014: data_o = 32'h00000000 /* 0x9c78 */;
                10015: data_o = 32'h00000000 /* 0x9c7c */;
                10016: data_o = 32'h00000000 /* 0x9c80 */;
                10017: data_o = 32'h00000000 /* 0x9c84 */;
                10018: data_o = 32'h00000000 /* 0x9c88 */;
                10019: data_o = 32'h00000000 /* 0x9c8c */;
                10020: data_o = 32'h00000000 /* 0x9c90 */;
                10021: data_o = 32'h00000000 /* 0x9c94 */;
                10022: data_o = 32'h00000000 /* 0x9c98 */;
                10023: data_o = 32'h00000000 /* 0x9c9c */;
                10024: data_o = 32'h00000000 /* 0x9ca0 */;
                10025: data_o = 32'h00000000 /* 0x9ca4 */;
                10026: data_o = 32'h00000000 /* 0x9ca8 */;
                10027: data_o = 32'h00000000 /* 0x9cac */;
                10028: data_o = 32'h00000000 /* 0x9cb0 */;
                10029: data_o = 32'h00000000 /* 0x9cb4 */;
                10030: data_o = 32'h00000000 /* 0x9cb8 */;
                10031: data_o = 32'h00000000 /* 0x9cbc */;
                10032: data_o = 32'h00000000 /* 0x9cc0 */;
                10033: data_o = 32'h00000000 /* 0x9cc4 */;
                10034: data_o = 32'h00000000 /* 0x9cc8 */;
                10035: data_o = 32'h00000000 /* 0x9ccc */;
                10036: data_o = 32'h00000000 /* 0x9cd0 */;
                10037: data_o = 32'h00000000 /* 0x9cd4 */;
                10038: data_o = 32'h00000000 /* 0x9cd8 */;
                10039: data_o = 32'h00000000 /* 0x9cdc */;
                10040: data_o = 32'h00000000 /* 0x9ce0 */;
                10041: data_o = 32'h00000000 /* 0x9ce4 */;
                10042: data_o = 32'h00000000 /* 0x9ce8 */;
                10043: data_o = 32'h00000000 /* 0x9cec */;
                10044: data_o = 32'h00000000 /* 0x9cf0 */;
                10045: data_o = 32'h00000000 /* 0x9cf4 */;
                10046: data_o = 32'h00000000 /* 0x9cf8 */;
                10047: data_o = 32'h00000000 /* 0x9cfc */;
                10048: data_o = 32'h00000000 /* 0x9d00 */;
                10049: data_o = 32'h00000000 /* 0x9d04 */;
                10050: data_o = 32'h00000000 /* 0x9d08 */;
                10051: data_o = 32'h00000000 /* 0x9d0c */;
                10052: data_o = 32'h00000000 /* 0x9d10 */;
                10053: data_o = 32'h00000000 /* 0x9d14 */;
                10054: data_o = 32'h00000000 /* 0x9d18 */;
                10055: data_o = 32'h00000000 /* 0x9d1c */;
                10056: data_o = 32'h00000000 /* 0x9d20 */;
                10057: data_o = 32'h00000000 /* 0x9d24 */;
                10058: data_o = 32'h00000000 /* 0x9d28 */;
                10059: data_o = 32'h00000000 /* 0x9d2c */;
                10060: data_o = 32'h00000000 /* 0x9d30 */;
                10061: data_o = 32'h00000000 /* 0x9d34 */;
                10062: data_o = 32'h00000000 /* 0x9d38 */;
                10063: data_o = 32'h00000000 /* 0x9d3c */;
                10064: data_o = 32'h00000000 /* 0x9d40 */;
                10065: data_o = 32'h00000000 /* 0x9d44 */;
                10066: data_o = 32'h00000000 /* 0x9d48 */;
                10067: data_o = 32'h00000000 /* 0x9d4c */;
                10068: data_o = 32'h00000000 /* 0x9d50 */;
                10069: data_o = 32'h00000000 /* 0x9d54 */;
                10070: data_o = 32'h00000000 /* 0x9d58 */;
                10071: data_o = 32'h00000000 /* 0x9d5c */;
                10072: data_o = 32'h00000000 /* 0x9d60 */;
                10073: data_o = 32'h00000000 /* 0x9d64 */;
                10074: data_o = 32'h00000000 /* 0x9d68 */;
                10075: data_o = 32'h00000000 /* 0x9d6c */;
                10076: data_o = 32'h00000000 /* 0x9d70 */;
                10077: data_o = 32'h00000000 /* 0x9d74 */;
                10078: data_o = 32'h00000000 /* 0x9d78 */;
                10079: data_o = 32'h00000000 /* 0x9d7c */;
                10080: data_o = 32'h00000000 /* 0x9d80 */;
                10081: data_o = 32'h00000000 /* 0x9d84 */;
                10082: data_o = 32'h00000000 /* 0x9d88 */;
                10083: data_o = 32'h00000000 /* 0x9d8c */;
                10084: data_o = 32'h00000000 /* 0x9d90 */;
                10085: data_o = 32'h00000000 /* 0x9d94 */;
                10086: data_o = 32'h00000000 /* 0x9d98 */;
                10087: data_o = 32'h00000000 /* 0x9d9c */;
                10088: data_o = 32'h00000000 /* 0x9da0 */;
                10089: data_o = 32'h00000000 /* 0x9da4 */;
                10090: data_o = 32'h00000000 /* 0x9da8 */;
                10091: data_o = 32'h00000000 /* 0x9dac */;
                10092: data_o = 32'h00000000 /* 0x9db0 */;
                10093: data_o = 32'h00000000 /* 0x9db4 */;
                10094: data_o = 32'h00000000 /* 0x9db8 */;
                10095: data_o = 32'h00000000 /* 0x9dbc */;
                10096: data_o = 32'h00000000 /* 0x9dc0 */;
                10097: data_o = 32'h00000000 /* 0x9dc4 */;
                10098: data_o = 32'h00000000 /* 0x9dc8 */;
                10099: data_o = 32'h00000000 /* 0x9dcc */;
                10100: data_o = 32'h00000000 /* 0x9dd0 */;
                10101: data_o = 32'h00000000 /* 0x9dd4 */;
                10102: data_o = 32'h00000000 /* 0x9dd8 */;
                10103: data_o = 32'h00000000 /* 0x9ddc */;
                10104: data_o = 32'h00000000 /* 0x9de0 */;
                10105: data_o = 32'h00000000 /* 0x9de4 */;
                10106: data_o = 32'h00000000 /* 0x9de8 */;
                10107: data_o = 32'h00000000 /* 0x9dec */;
                10108: data_o = 32'h00000000 /* 0x9df0 */;
                10109: data_o = 32'h00000000 /* 0x9df4 */;
                10110: data_o = 32'h00000000 /* 0x9df8 */;
                10111: data_o = 32'h00000000 /* 0x9dfc */;
                10112: data_o = 32'h00000000 /* 0x9e00 */;
                10113: data_o = 32'h00000000 /* 0x9e04 */;
                10114: data_o = 32'h00000000 /* 0x9e08 */;
                10115: data_o = 32'h00000000 /* 0x9e0c */;
                10116: data_o = 32'h00000000 /* 0x9e10 */;
                10117: data_o = 32'h00000000 /* 0x9e14 */;
                10118: data_o = 32'h00000000 /* 0x9e18 */;
                10119: data_o = 32'h00000000 /* 0x9e1c */;
                10120: data_o = 32'h00000000 /* 0x9e20 */;
                10121: data_o = 32'h00000000 /* 0x9e24 */;
                10122: data_o = 32'h00000000 /* 0x9e28 */;
                10123: data_o = 32'h00000000 /* 0x9e2c */;
                10124: data_o = 32'h00000000 /* 0x9e30 */;
                10125: data_o = 32'h00000000 /* 0x9e34 */;
                10126: data_o = 32'h00000000 /* 0x9e38 */;
                10127: data_o = 32'h00000000 /* 0x9e3c */;
                10128: data_o = 32'h00000000 /* 0x9e40 */;
                10129: data_o = 32'h00000000 /* 0x9e44 */;
                10130: data_o = 32'h00000000 /* 0x9e48 */;
                10131: data_o = 32'h00000000 /* 0x9e4c */;
                10132: data_o = 32'h00000000 /* 0x9e50 */;
                10133: data_o = 32'h00000000 /* 0x9e54 */;
                10134: data_o = 32'h00000000 /* 0x9e58 */;
                10135: data_o = 32'h00000000 /* 0x9e5c */;
                10136: data_o = 32'h00000000 /* 0x9e60 */;
                10137: data_o = 32'h00000000 /* 0x9e64 */;
                10138: data_o = 32'h00000000 /* 0x9e68 */;
                10139: data_o = 32'h00000000 /* 0x9e6c */;
                10140: data_o = 32'h00000000 /* 0x9e70 */;
                10141: data_o = 32'h00000000 /* 0x9e74 */;
                10142: data_o = 32'h00000000 /* 0x9e78 */;
                10143: data_o = 32'h00000000 /* 0x9e7c */;
                10144: data_o = 32'h00000000 /* 0x9e80 */;
                10145: data_o = 32'h00000000 /* 0x9e84 */;
                10146: data_o = 32'h00000000 /* 0x9e88 */;
                10147: data_o = 32'h00000000 /* 0x9e8c */;
                10148: data_o = 32'h00000000 /* 0x9e90 */;
                10149: data_o = 32'h00000000 /* 0x9e94 */;
                10150: data_o = 32'h00000000 /* 0x9e98 */;
                10151: data_o = 32'h00000000 /* 0x9e9c */;
                10152: data_o = 32'h00000000 /* 0x9ea0 */;
                10153: data_o = 32'h00000000 /* 0x9ea4 */;
                10154: data_o = 32'h00000000 /* 0x9ea8 */;
                10155: data_o = 32'h00000000 /* 0x9eac */;
                10156: data_o = 32'h00000000 /* 0x9eb0 */;
                10157: data_o = 32'h00000000 /* 0x9eb4 */;
                10158: data_o = 32'h00000000 /* 0x9eb8 */;
                10159: data_o = 32'h00000000 /* 0x9ebc */;
                10160: data_o = 32'h00000000 /* 0x9ec0 */;
                10161: data_o = 32'h00000000 /* 0x9ec4 */;
                10162: data_o = 32'h00000000 /* 0x9ec8 */;
                10163: data_o = 32'h00000000 /* 0x9ecc */;
                10164: data_o = 32'h00000000 /* 0x9ed0 */;
                10165: data_o = 32'h00000000 /* 0x9ed4 */;
                10166: data_o = 32'h00000000 /* 0x9ed8 */;
                10167: data_o = 32'h00000000 /* 0x9edc */;
                10168: data_o = 32'h00000000 /* 0x9ee0 */;
                10169: data_o = 32'h00000000 /* 0x9ee4 */;
                10170: data_o = 32'h00000000 /* 0x9ee8 */;
                10171: data_o = 32'h00000000 /* 0x9eec */;
                10172: data_o = 32'h00000000 /* 0x9ef0 */;
                10173: data_o = 32'h00000000 /* 0x9ef4 */;
                10174: data_o = 32'h00000000 /* 0x9ef8 */;
                10175: data_o = 32'h00000000 /* 0x9efc */;
                10176: data_o = 32'h00000000 /* 0x9f00 */;
                10177: data_o = 32'h00000000 /* 0x9f04 */;
                10178: data_o = 32'h00000000 /* 0x9f08 */;
                10179: data_o = 32'h00000000 /* 0x9f0c */;
                10180: data_o = 32'h00000000 /* 0x9f10 */;
                10181: data_o = 32'h00000000 /* 0x9f14 */;
                10182: data_o = 32'h00000000 /* 0x9f18 */;
                10183: data_o = 32'h00000000 /* 0x9f1c */;
                10184: data_o = 32'h00000000 /* 0x9f20 */;
                10185: data_o = 32'h00000000 /* 0x9f24 */;
                10186: data_o = 32'h00000000 /* 0x9f28 */;
                10187: data_o = 32'h00000000 /* 0x9f2c */;
                10188: data_o = 32'h00000000 /* 0x9f30 */;
                10189: data_o = 32'h00000000 /* 0x9f34 */;
                10190: data_o = 32'h00000000 /* 0x9f38 */;
                10191: data_o = 32'h00000000 /* 0x9f3c */;
                10192: data_o = 32'h00000000 /* 0x9f40 */;
                10193: data_o = 32'h00000000 /* 0x9f44 */;
                10194: data_o = 32'h00000000 /* 0x9f48 */;
                10195: data_o = 32'h00000000 /* 0x9f4c */;
                10196: data_o = 32'h00000000 /* 0x9f50 */;
                10197: data_o = 32'h00000000 /* 0x9f54 */;
                10198: data_o = 32'h00000000 /* 0x9f58 */;
                10199: data_o = 32'h00000000 /* 0x9f5c */;
                10200: data_o = 32'h00000000 /* 0x9f60 */;
                10201: data_o = 32'h00000000 /* 0x9f64 */;
                10202: data_o = 32'h00000000 /* 0x9f68 */;
                10203: data_o = 32'h00000000 /* 0x9f6c */;
                10204: data_o = 32'h00000000 /* 0x9f70 */;
                10205: data_o = 32'h00000000 /* 0x9f74 */;
                10206: data_o = 32'h00000000 /* 0x9f78 */;
                10207: data_o = 32'h00000000 /* 0x9f7c */;
                10208: data_o = 32'h00000000 /* 0x9f80 */;
                10209: data_o = 32'h00000000 /* 0x9f84 */;
                10210: data_o = 32'h00000000 /* 0x9f88 */;
                10211: data_o = 32'h00000000 /* 0x9f8c */;
                10212: data_o = 32'h00000000 /* 0x9f90 */;
                10213: data_o = 32'h00000000 /* 0x9f94 */;
                10214: data_o = 32'h00000000 /* 0x9f98 */;
                10215: data_o = 32'h00000000 /* 0x9f9c */;
                10216: data_o = 32'h00000000 /* 0x9fa0 */;
                10217: data_o = 32'h00000000 /* 0x9fa4 */;
                10218: data_o = 32'h00000000 /* 0x9fa8 */;
                10219: data_o = 32'h00000000 /* 0x9fac */;
                10220: data_o = 32'h00000000 /* 0x9fb0 */;
                10221: data_o = 32'h00000000 /* 0x9fb4 */;
                10222: data_o = 32'h00000000 /* 0x9fb8 */;
                10223: data_o = 32'h00000000 /* 0x9fbc */;
                10224: data_o = 32'h00000000 /* 0x9fc0 */;
                10225: data_o = 32'h00000000 /* 0x9fc4 */;
                10226: data_o = 32'h00000000 /* 0x9fc8 */;
                10227: data_o = 32'h00000000 /* 0x9fcc */;
                10228: data_o = 32'h00000000 /* 0x9fd0 */;
                10229: data_o = 32'h00000000 /* 0x9fd4 */;
                10230: data_o = 32'h00000000 /* 0x9fd8 */;
                10231: data_o = 32'h00000000 /* 0x9fdc */;
                10232: data_o = 32'h00000000 /* 0x9fe0 */;
                10233: data_o = 32'h00000000 /* 0x9fe4 */;
                10234: data_o = 32'h00000000 /* 0x9fe8 */;
                10235: data_o = 32'h00000000 /* 0x9fec */;
                10236: data_o = 32'h00000000 /* 0x9ff0 */;
                10237: data_o = 32'h00000000 /* 0x9ff4 */;
                10238: data_o = 32'h00000000 /* 0x9ff8 */;
                10239: data_o = 32'h00000000 /* 0x9ffc */;
                10240: data_o = 32'h00000000 /* 0xa000 */;
                10241: data_o = 32'h00000000 /* 0xa004 */;
                10242: data_o = 32'h00000000 /* 0xa008 */;
                10243: data_o = 32'h00000000 /* 0xa00c */;
                10244: data_o = 32'h00000000 /* 0xa010 */;
                10245: data_o = 32'h00000000 /* 0xa014 */;
                10246: data_o = 32'h00000000 /* 0xa018 */;
                10247: data_o = 32'h00000000 /* 0xa01c */;
                10248: data_o = 32'h00000000 /* 0xa020 */;
                10249: data_o = 32'h00000000 /* 0xa024 */;
                10250: data_o = 32'h00000000 /* 0xa028 */;
                10251: data_o = 32'h00000000 /* 0xa02c */;
                10252: data_o = 32'h00000000 /* 0xa030 */;
                10253: data_o = 32'h00000000 /* 0xa034 */;
                10254: data_o = 32'h00000000 /* 0xa038 */;
                10255: data_o = 32'h00000000 /* 0xa03c */;
                10256: data_o = 32'h00000000 /* 0xa040 */;
                10257: data_o = 32'h00000000 /* 0xa044 */;
                10258: data_o = 32'h00000000 /* 0xa048 */;
                10259: data_o = 32'h00000000 /* 0xa04c */;
                10260: data_o = 32'h00000000 /* 0xa050 */;
                10261: data_o = 32'h00000000 /* 0xa054 */;
                10262: data_o = 32'h00000000 /* 0xa058 */;
                10263: data_o = 32'h00000000 /* 0xa05c */;
                10264: data_o = 32'h00000000 /* 0xa060 */;
                10265: data_o = 32'h00000000 /* 0xa064 */;
                10266: data_o = 32'h00000000 /* 0xa068 */;
                10267: data_o = 32'h00000000 /* 0xa06c */;
                10268: data_o = 32'h00000000 /* 0xa070 */;
                10269: data_o = 32'h00000000 /* 0xa074 */;
                10270: data_o = 32'h00000000 /* 0xa078 */;
                10271: data_o = 32'h00000000 /* 0xa07c */;
                10272: data_o = 32'h00000000 /* 0xa080 */;
                10273: data_o = 32'h00000000 /* 0xa084 */;
                10274: data_o = 32'h00000000 /* 0xa088 */;
                10275: data_o = 32'h00000000 /* 0xa08c */;
                10276: data_o = 32'h00000000 /* 0xa090 */;
                10277: data_o = 32'h00000000 /* 0xa094 */;
                10278: data_o = 32'h00000000 /* 0xa098 */;
                10279: data_o = 32'h00000000 /* 0xa09c */;
                10280: data_o = 32'h00000000 /* 0xa0a0 */;
                10281: data_o = 32'h00000000 /* 0xa0a4 */;
                10282: data_o = 32'h00000000 /* 0xa0a8 */;
                10283: data_o = 32'h00000000 /* 0xa0ac */;
                10284: data_o = 32'h00000000 /* 0xa0b0 */;
                10285: data_o = 32'h00000000 /* 0xa0b4 */;
                10286: data_o = 32'h00000000 /* 0xa0b8 */;
                10287: data_o = 32'h00000000 /* 0xa0bc */;
                10288: data_o = 32'h00000000 /* 0xa0c0 */;
                10289: data_o = 32'h00000000 /* 0xa0c4 */;
                10290: data_o = 32'h00000000 /* 0xa0c8 */;
                10291: data_o = 32'h00000000 /* 0xa0cc */;
                10292: data_o = 32'h00000000 /* 0xa0d0 */;
                10293: data_o = 32'h00000000 /* 0xa0d4 */;
                10294: data_o = 32'h00000000 /* 0xa0d8 */;
                10295: data_o = 32'h00000000 /* 0xa0dc */;
                10296: data_o = 32'h00000000 /* 0xa0e0 */;
                10297: data_o = 32'h00000000 /* 0xa0e4 */;
                10298: data_o = 32'h00000000 /* 0xa0e8 */;
                10299: data_o = 32'h00000000 /* 0xa0ec */;
                10300: data_o = 32'h00000000 /* 0xa0f0 */;
                10301: data_o = 32'h00000000 /* 0xa0f4 */;
                10302: data_o = 32'h00000000 /* 0xa0f8 */;
                10303: data_o = 32'h00000000 /* 0xa0fc */;
                10304: data_o = 32'h00000000 /* 0xa100 */;
                10305: data_o = 32'h00000000 /* 0xa104 */;
                10306: data_o = 32'h00000000 /* 0xa108 */;
                10307: data_o = 32'h00000000 /* 0xa10c */;
                10308: data_o = 32'h00000000 /* 0xa110 */;
                10309: data_o = 32'h00000000 /* 0xa114 */;
                10310: data_o = 32'h00000000 /* 0xa118 */;
                10311: data_o = 32'h00000000 /* 0xa11c */;
                10312: data_o = 32'h00000000 /* 0xa120 */;
                10313: data_o = 32'h00000000 /* 0xa124 */;
                10314: data_o = 32'h00000000 /* 0xa128 */;
                10315: data_o = 32'h00000000 /* 0xa12c */;
                10316: data_o = 32'h00000000 /* 0xa130 */;
                10317: data_o = 32'h00000000 /* 0xa134 */;
                10318: data_o = 32'h00000000 /* 0xa138 */;
                10319: data_o = 32'h00000000 /* 0xa13c */;
                10320: data_o = 32'h00000000 /* 0xa140 */;
                10321: data_o = 32'h00000000 /* 0xa144 */;
                10322: data_o = 32'h00000000 /* 0xa148 */;
                10323: data_o = 32'h00000000 /* 0xa14c */;
                10324: data_o = 32'h00000000 /* 0xa150 */;
                10325: data_o = 32'h00000000 /* 0xa154 */;
                10326: data_o = 32'h00000000 /* 0xa158 */;
                10327: data_o = 32'h00000000 /* 0xa15c */;
                10328: data_o = 32'h00000000 /* 0xa160 */;
                10329: data_o = 32'h00000000 /* 0xa164 */;
                10330: data_o = 32'h00000000 /* 0xa168 */;
                10331: data_o = 32'h00000000 /* 0xa16c */;
                10332: data_o = 32'h00000000 /* 0xa170 */;
                10333: data_o = 32'h00000000 /* 0xa174 */;
                10334: data_o = 32'h00000000 /* 0xa178 */;
                10335: data_o = 32'h00000000 /* 0xa17c */;
                10336: data_o = 32'h00000000 /* 0xa180 */;
                10337: data_o = 32'h00000000 /* 0xa184 */;
                10338: data_o = 32'h00000000 /* 0xa188 */;
                10339: data_o = 32'h00000000 /* 0xa18c */;
                10340: data_o = 32'h00000000 /* 0xa190 */;
                10341: data_o = 32'h00000000 /* 0xa194 */;
                10342: data_o = 32'h00000000 /* 0xa198 */;
                10343: data_o = 32'h00000000 /* 0xa19c */;
                10344: data_o = 32'h00000000 /* 0xa1a0 */;
                10345: data_o = 32'h00000000 /* 0xa1a4 */;
                10346: data_o = 32'h00000000 /* 0xa1a8 */;
                10347: data_o = 32'h00000000 /* 0xa1ac */;
                10348: data_o = 32'h00000000 /* 0xa1b0 */;
                10349: data_o = 32'h00000000 /* 0xa1b4 */;
                10350: data_o = 32'h00000000 /* 0xa1b8 */;
                10351: data_o = 32'h00000000 /* 0xa1bc */;
                10352: data_o = 32'h00000000 /* 0xa1c0 */;
                10353: data_o = 32'h00000000 /* 0xa1c4 */;
                10354: data_o = 32'h00000000 /* 0xa1c8 */;
                10355: data_o = 32'h00000000 /* 0xa1cc */;
                10356: data_o = 32'h00000000 /* 0xa1d0 */;
                10357: data_o = 32'h00000000 /* 0xa1d4 */;
                10358: data_o = 32'h00000000 /* 0xa1d8 */;
                10359: data_o = 32'h00000000 /* 0xa1dc */;
                10360: data_o = 32'h00000000 /* 0xa1e0 */;
                10361: data_o = 32'h00000000 /* 0xa1e4 */;
                10362: data_o = 32'h00000000 /* 0xa1e8 */;
                10363: data_o = 32'h00000000 /* 0xa1ec */;
                10364: data_o = 32'h00000000 /* 0xa1f0 */;
                10365: data_o = 32'h00000000 /* 0xa1f4 */;
                10366: data_o = 32'h00000000 /* 0xa1f8 */;
                10367: data_o = 32'h00000000 /* 0xa1fc */;
                10368: data_o = 32'h00000000 /* 0xa200 */;
                10369: data_o = 32'h00000000 /* 0xa204 */;
                10370: data_o = 32'h00000000 /* 0xa208 */;
                10371: data_o = 32'h00000000 /* 0xa20c */;
                10372: data_o = 32'h00000000 /* 0xa210 */;
                10373: data_o = 32'h00000000 /* 0xa214 */;
                10374: data_o = 32'h00000000 /* 0xa218 */;
                10375: data_o = 32'h00000000 /* 0xa21c */;
                10376: data_o = 32'h00000000 /* 0xa220 */;
                10377: data_o = 32'h00000000 /* 0xa224 */;
                10378: data_o = 32'h00000000 /* 0xa228 */;
                10379: data_o = 32'h00000000 /* 0xa22c */;
                10380: data_o = 32'h00000000 /* 0xa230 */;
                10381: data_o = 32'h00000000 /* 0xa234 */;
                10382: data_o = 32'h00000000 /* 0xa238 */;
                10383: data_o = 32'h00000000 /* 0xa23c */;
                10384: data_o = 32'h00000000 /* 0xa240 */;
                10385: data_o = 32'h00000000 /* 0xa244 */;
                10386: data_o = 32'h00000000 /* 0xa248 */;
                10387: data_o = 32'h00000000 /* 0xa24c */;
                10388: data_o = 32'h00000000 /* 0xa250 */;
                10389: data_o = 32'h00000000 /* 0xa254 */;
                10390: data_o = 32'h00000000 /* 0xa258 */;
                10391: data_o = 32'h00000000 /* 0xa25c */;
                10392: data_o = 32'h00000000 /* 0xa260 */;
                10393: data_o = 32'h00000000 /* 0xa264 */;
                10394: data_o = 32'h00000000 /* 0xa268 */;
                10395: data_o = 32'h00000000 /* 0xa26c */;
                10396: data_o = 32'h00000000 /* 0xa270 */;
                10397: data_o = 32'h00000000 /* 0xa274 */;
                10398: data_o = 32'h00000000 /* 0xa278 */;
                10399: data_o = 32'h00000000 /* 0xa27c */;
                10400: data_o = 32'h00000000 /* 0xa280 */;
                10401: data_o = 32'h00000000 /* 0xa284 */;
                10402: data_o = 32'h00000000 /* 0xa288 */;
                10403: data_o = 32'h00000000 /* 0xa28c */;
                10404: data_o = 32'h00000000 /* 0xa290 */;
                10405: data_o = 32'h00000000 /* 0xa294 */;
                10406: data_o = 32'h00000000 /* 0xa298 */;
                10407: data_o = 32'h00000000 /* 0xa29c */;
                10408: data_o = 32'h00000000 /* 0xa2a0 */;
                10409: data_o = 32'h00000000 /* 0xa2a4 */;
                10410: data_o = 32'h00000000 /* 0xa2a8 */;
                10411: data_o = 32'h00000000 /* 0xa2ac */;
                10412: data_o = 32'h00000000 /* 0xa2b0 */;
                10413: data_o = 32'h00000000 /* 0xa2b4 */;
                10414: data_o = 32'h00000000 /* 0xa2b8 */;
                10415: data_o = 32'h00000000 /* 0xa2bc */;
                10416: data_o = 32'h00000000 /* 0xa2c0 */;
                10417: data_o = 32'h00000000 /* 0xa2c4 */;
                10418: data_o = 32'h00000000 /* 0xa2c8 */;
                10419: data_o = 32'h00000000 /* 0xa2cc */;
                10420: data_o = 32'h00000000 /* 0xa2d0 */;
                10421: data_o = 32'h00000000 /* 0xa2d4 */;
                10422: data_o = 32'h00000000 /* 0xa2d8 */;
                10423: data_o = 32'h00000000 /* 0xa2dc */;
                10424: data_o = 32'h00000000 /* 0xa2e0 */;
                10425: data_o = 32'h00000000 /* 0xa2e4 */;
                10426: data_o = 32'h00000000 /* 0xa2e8 */;
                10427: data_o = 32'h00000000 /* 0xa2ec */;
                10428: data_o = 32'h00000000 /* 0xa2f0 */;
                10429: data_o = 32'h00000000 /* 0xa2f4 */;
                10430: data_o = 32'h00000000 /* 0xa2f8 */;
                10431: data_o = 32'h00000000 /* 0xa2fc */;
                10432: data_o = 32'h00000000 /* 0xa300 */;
                10433: data_o = 32'h00000000 /* 0xa304 */;
                10434: data_o = 32'h00000000 /* 0xa308 */;
                10435: data_o = 32'h00000000 /* 0xa30c */;
                10436: data_o = 32'h00000000 /* 0xa310 */;
                10437: data_o = 32'h00000000 /* 0xa314 */;
                10438: data_o = 32'h00000000 /* 0xa318 */;
                10439: data_o = 32'h00000000 /* 0xa31c */;
                10440: data_o = 32'h00000000 /* 0xa320 */;
                10441: data_o = 32'h00000000 /* 0xa324 */;
                10442: data_o = 32'h00000000 /* 0xa328 */;
                10443: data_o = 32'h00000000 /* 0xa32c */;
                10444: data_o = 32'h00000000 /* 0xa330 */;
                10445: data_o = 32'h00000000 /* 0xa334 */;
                10446: data_o = 32'h00000000 /* 0xa338 */;
                10447: data_o = 32'h00000000 /* 0xa33c */;
                10448: data_o = 32'h00000000 /* 0xa340 */;
                10449: data_o = 32'h00000000 /* 0xa344 */;
                10450: data_o = 32'h00000000 /* 0xa348 */;
                10451: data_o = 32'h00000000 /* 0xa34c */;
                10452: data_o = 32'h00000000 /* 0xa350 */;
                10453: data_o = 32'h00000000 /* 0xa354 */;
                10454: data_o = 32'h00000000 /* 0xa358 */;
                10455: data_o = 32'h00000000 /* 0xa35c */;
                10456: data_o = 32'h00000000 /* 0xa360 */;
                10457: data_o = 32'h00000000 /* 0xa364 */;
                10458: data_o = 32'h00000000 /* 0xa368 */;
                10459: data_o = 32'h00000000 /* 0xa36c */;
                10460: data_o = 32'h00000000 /* 0xa370 */;
                10461: data_o = 32'h00000000 /* 0xa374 */;
                10462: data_o = 32'h00000000 /* 0xa378 */;
                10463: data_o = 32'h00000000 /* 0xa37c */;
                10464: data_o = 32'h00000000 /* 0xa380 */;
                10465: data_o = 32'h00000000 /* 0xa384 */;
                10466: data_o = 32'h00000000 /* 0xa388 */;
                10467: data_o = 32'h00000000 /* 0xa38c */;
                10468: data_o = 32'h00000000 /* 0xa390 */;
                10469: data_o = 32'h00000000 /* 0xa394 */;
                10470: data_o = 32'h00000000 /* 0xa398 */;
                10471: data_o = 32'h00000000 /* 0xa39c */;
                10472: data_o = 32'h00000000 /* 0xa3a0 */;
                10473: data_o = 32'h00000000 /* 0xa3a4 */;
                10474: data_o = 32'h00000000 /* 0xa3a8 */;
                10475: data_o = 32'h00000000 /* 0xa3ac */;
                10476: data_o = 32'h00000000 /* 0xa3b0 */;
                10477: data_o = 32'h00000000 /* 0xa3b4 */;
                10478: data_o = 32'h00000000 /* 0xa3b8 */;
                10479: data_o = 32'h00000000 /* 0xa3bc */;
                10480: data_o = 32'h00000000 /* 0xa3c0 */;
                10481: data_o = 32'h00000000 /* 0xa3c4 */;
                10482: data_o = 32'h00000000 /* 0xa3c8 */;
                10483: data_o = 32'h00000000 /* 0xa3cc */;
                10484: data_o = 32'h00000000 /* 0xa3d0 */;
                10485: data_o = 32'h00000000 /* 0xa3d4 */;
                10486: data_o = 32'h00000000 /* 0xa3d8 */;
                10487: data_o = 32'h00000000 /* 0xa3dc */;
                10488: data_o = 32'h00000000 /* 0xa3e0 */;
                10489: data_o = 32'h00000000 /* 0xa3e4 */;
                10490: data_o = 32'h00000000 /* 0xa3e8 */;
                10491: data_o = 32'h00000000 /* 0xa3ec */;
                10492: data_o = 32'h00000000 /* 0xa3f0 */;
                10493: data_o = 32'h00000000 /* 0xa3f4 */;
                10494: data_o = 32'h00000000 /* 0xa3f8 */;
                10495: data_o = 32'h00000000 /* 0xa3fc */;
                10496: data_o = 32'h00000000 /* 0xa400 */;
                10497: data_o = 32'h00000000 /* 0xa404 */;
                10498: data_o = 32'h00000000 /* 0xa408 */;
                10499: data_o = 32'h00000000 /* 0xa40c */;
                10500: data_o = 32'h00000000 /* 0xa410 */;
                10501: data_o = 32'h00000000 /* 0xa414 */;
                10502: data_o = 32'h00000000 /* 0xa418 */;
                10503: data_o = 32'h00000000 /* 0xa41c */;
                10504: data_o = 32'h00000000 /* 0xa420 */;
                10505: data_o = 32'h00000000 /* 0xa424 */;
                10506: data_o = 32'h00000000 /* 0xa428 */;
                10507: data_o = 32'h00000000 /* 0xa42c */;
                10508: data_o = 32'h00000000 /* 0xa430 */;
                10509: data_o = 32'h00000000 /* 0xa434 */;
                10510: data_o = 32'h00000000 /* 0xa438 */;
                10511: data_o = 32'h00000000 /* 0xa43c */;
                10512: data_o = 32'h00000000 /* 0xa440 */;
                10513: data_o = 32'h00000000 /* 0xa444 */;
                10514: data_o = 32'h00000000 /* 0xa448 */;
                10515: data_o = 32'h00000000 /* 0xa44c */;
                10516: data_o = 32'h00000000 /* 0xa450 */;
                10517: data_o = 32'h00000000 /* 0xa454 */;
                10518: data_o = 32'h00000000 /* 0xa458 */;
                10519: data_o = 32'h00000000 /* 0xa45c */;
                10520: data_o = 32'h00000000 /* 0xa460 */;
                10521: data_o = 32'h00000000 /* 0xa464 */;
                10522: data_o = 32'h00000000 /* 0xa468 */;
                10523: data_o = 32'h00000000 /* 0xa46c */;
                10524: data_o = 32'h00000000 /* 0xa470 */;
                10525: data_o = 32'h00000000 /* 0xa474 */;
                10526: data_o = 32'h00000000 /* 0xa478 */;
                10527: data_o = 32'h00000000 /* 0xa47c */;
                10528: data_o = 32'h00000000 /* 0xa480 */;
                10529: data_o = 32'h00000000 /* 0xa484 */;
                10530: data_o = 32'h00000000 /* 0xa488 */;
                10531: data_o = 32'h00000000 /* 0xa48c */;
                10532: data_o = 32'h00000000 /* 0xa490 */;
                10533: data_o = 32'h00000000 /* 0xa494 */;
                10534: data_o = 32'h00000000 /* 0xa498 */;
                10535: data_o = 32'h00000000 /* 0xa49c */;
                10536: data_o = 32'h00000000 /* 0xa4a0 */;
                10537: data_o = 32'h00000000 /* 0xa4a4 */;
                10538: data_o = 32'h00000000 /* 0xa4a8 */;
                10539: data_o = 32'h00000000 /* 0xa4ac */;
                10540: data_o = 32'h00000000 /* 0xa4b0 */;
                10541: data_o = 32'h00000000 /* 0xa4b4 */;
                10542: data_o = 32'h00000000 /* 0xa4b8 */;
                10543: data_o = 32'h00000000 /* 0xa4bc */;
                10544: data_o = 32'h00000000 /* 0xa4c0 */;
                10545: data_o = 32'h00000000 /* 0xa4c4 */;
                10546: data_o = 32'h00000000 /* 0xa4c8 */;
                10547: data_o = 32'h00000000 /* 0xa4cc */;
                10548: data_o = 32'h00000000 /* 0xa4d0 */;
                10549: data_o = 32'h00000000 /* 0xa4d4 */;
                10550: data_o = 32'h00000000 /* 0xa4d8 */;
                10551: data_o = 32'h00000000 /* 0xa4dc */;
                10552: data_o = 32'h00000000 /* 0xa4e0 */;
                10553: data_o = 32'h00000000 /* 0xa4e4 */;
                10554: data_o = 32'h00000000 /* 0xa4e8 */;
                10555: data_o = 32'h00000000 /* 0xa4ec */;
                10556: data_o = 32'h00000000 /* 0xa4f0 */;
                10557: data_o = 32'h00000000 /* 0xa4f4 */;
                10558: data_o = 32'h00000000 /* 0xa4f8 */;
                10559: data_o = 32'h00000000 /* 0xa4fc */;
                10560: data_o = 32'h00000000 /* 0xa500 */;
                10561: data_o = 32'h00000000 /* 0xa504 */;
                10562: data_o = 32'h00000000 /* 0xa508 */;
                10563: data_o = 32'h00000000 /* 0xa50c */;
                10564: data_o = 32'h00000000 /* 0xa510 */;
                10565: data_o = 32'h00000000 /* 0xa514 */;
                10566: data_o = 32'h00000000 /* 0xa518 */;
                10567: data_o = 32'h00000000 /* 0xa51c */;
                10568: data_o = 32'h00000000 /* 0xa520 */;
                10569: data_o = 32'h00000000 /* 0xa524 */;
                10570: data_o = 32'h00000000 /* 0xa528 */;
                10571: data_o = 32'h00000000 /* 0xa52c */;
                10572: data_o = 32'h00000000 /* 0xa530 */;
                10573: data_o = 32'h00000000 /* 0xa534 */;
                10574: data_o = 32'h00000000 /* 0xa538 */;
                10575: data_o = 32'h00000000 /* 0xa53c */;
                10576: data_o = 32'h00000000 /* 0xa540 */;
                10577: data_o = 32'h00000000 /* 0xa544 */;
                10578: data_o = 32'h00000000 /* 0xa548 */;
                10579: data_o = 32'h00000000 /* 0xa54c */;
                10580: data_o = 32'h00000000 /* 0xa550 */;
                10581: data_o = 32'h00000000 /* 0xa554 */;
                10582: data_o = 32'h00000000 /* 0xa558 */;
                10583: data_o = 32'h00000000 /* 0xa55c */;
                10584: data_o = 32'h00000000 /* 0xa560 */;
                10585: data_o = 32'h00000000 /* 0xa564 */;
                10586: data_o = 32'h00000000 /* 0xa568 */;
                10587: data_o = 32'h00000000 /* 0xa56c */;
                10588: data_o = 32'h00000000 /* 0xa570 */;
                10589: data_o = 32'h00000000 /* 0xa574 */;
                10590: data_o = 32'h00000000 /* 0xa578 */;
                10591: data_o = 32'h00000000 /* 0xa57c */;
                10592: data_o = 32'h00000000 /* 0xa580 */;
                10593: data_o = 32'h00000000 /* 0xa584 */;
                10594: data_o = 32'h00000000 /* 0xa588 */;
                10595: data_o = 32'h00000000 /* 0xa58c */;
                10596: data_o = 32'h00000000 /* 0xa590 */;
                10597: data_o = 32'h00000000 /* 0xa594 */;
                10598: data_o = 32'h00000000 /* 0xa598 */;
                10599: data_o = 32'h00000000 /* 0xa59c */;
                10600: data_o = 32'h00000000 /* 0xa5a0 */;
                10601: data_o = 32'h00000000 /* 0xa5a4 */;
                10602: data_o = 32'h00000000 /* 0xa5a8 */;
                10603: data_o = 32'h00000000 /* 0xa5ac */;
                10604: data_o = 32'h00000000 /* 0xa5b0 */;
                10605: data_o = 32'h00000000 /* 0xa5b4 */;
                10606: data_o = 32'h00000000 /* 0xa5b8 */;
                10607: data_o = 32'h00000000 /* 0xa5bc */;
                10608: data_o = 32'h00000000 /* 0xa5c0 */;
                10609: data_o = 32'h00000000 /* 0xa5c4 */;
                10610: data_o = 32'h00000000 /* 0xa5c8 */;
                10611: data_o = 32'h00000000 /* 0xa5cc */;
                10612: data_o = 32'h00000000 /* 0xa5d0 */;
                10613: data_o = 32'h00000000 /* 0xa5d4 */;
                10614: data_o = 32'h00000000 /* 0xa5d8 */;
                10615: data_o = 32'h00000000 /* 0xa5dc */;
                10616: data_o = 32'h00000000 /* 0xa5e0 */;
                10617: data_o = 32'h00000000 /* 0xa5e4 */;
                10618: data_o = 32'h00000000 /* 0xa5e8 */;
                10619: data_o = 32'h00000000 /* 0xa5ec */;
                10620: data_o = 32'h00000000 /* 0xa5f0 */;
                10621: data_o = 32'h00000000 /* 0xa5f4 */;
                10622: data_o = 32'h00000000 /* 0xa5f8 */;
                10623: data_o = 32'h00000000 /* 0xa5fc */;
                10624: data_o = 32'h00000000 /* 0xa600 */;
                10625: data_o = 32'h00000000 /* 0xa604 */;
                10626: data_o = 32'h00000000 /* 0xa608 */;
                10627: data_o = 32'h00000000 /* 0xa60c */;
                10628: data_o = 32'h00000000 /* 0xa610 */;
                10629: data_o = 32'h00000000 /* 0xa614 */;
                10630: data_o = 32'h00000000 /* 0xa618 */;
                10631: data_o = 32'h00000000 /* 0xa61c */;
                10632: data_o = 32'h00000000 /* 0xa620 */;
                10633: data_o = 32'h00000000 /* 0xa624 */;
                10634: data_o = 32'h00000000 /* 0xa628 */;
                10635: data_o = 32'h00000000 /* 0xa62c */;
                10636: data_o = 32'h00000000 /* 0xa630 */;
                10637: data_o = 32'h00000000 /* 0xa634 */;
                10638: data_o = 32'h00000000 /* 0xa638 */;
                10639: data_o = 32'h00000000 /* 0xa63c */;
                10640: data_o = 32'h00000000 /* 0xa640 */;
                10641: data_o = 32'h00000000 /* 0xa644 */;
                10642: data_o = 32'h00000000 /* 0xa648 */;
                10643: data_o = 32'h00000000 /* 0xa64c */;
                10644: data_o = 32'h00000000 /* 0xa650 */;
                10645: data_o = 32'h00000000 /* 0xa654 */;
                10646: data_o = 32'h00000000 /* 0xa658 */;
                10647: data_o = 32'h00000000 /* 0xa65c */;
                10648: data_o = 32'h00000000 /* 0xa660 */;
                10649: data_o = 32'h00000000 /* 0xa664 */;
                10650: data_o = 32'h00000000 /* 0xa668 */;
                10651: data_o = 32'h00000000 /* 0xa66c */;
                10652: data_o = 32'h00000000 /* 0xa670 */;
                10653: data_o = 32'h00000000 /* 0xa674 */;
                10654: data_o = 32'h00000000 /* 0xa678 */;
                10655: data_o = 32'h00000000 /* 0xa67c */;
                10656: data_o = 32'h00000000 /* 0xa680 */;
                10657: data_o = 32'h00000000 /* 0xa684 */;
                10658: data_o = 32'h00000000 /* 0xa688 */;
                10659: data_o = 32'h00000000 /* 0xa68c */;
                10660: data_o = 32'h00000000 /* 0xa690 */;
                10661: data_o = 32'h00000000 /* 0xa694 */;
                10662: data_o = 32'h00000000 /* 0xa698 */;
                10663: data_o = 32'h00000000 /* 0xa69c */;
                10664: data_o = 32'h00000000 /* 0xa6a0 */;
                10665: data_o = 32'h00000000 /* 0xa6a4 */;
                10666: data_o = 32'h00000000 /* 0xa6a8 */;
                10667: data_o = 32'h00000000 /* 0xa6ac */;
                10668: data_o = 32'h00000000 /* 0xa6b0 */;
                10669: data_o = 32'h00000000 /* 0xa6b4 */;
                10670: data_o = 32'h00000000 /* 0xa6b8 */;
                10671: data_o = 32'h00000000 /* 0xa6bc */;
                10672: data_o = 32'h00000000 /* 0xa6c0 */;
                10673: data_o = 32'h00000000 /* 0xa6c4 */;
                10674: data_o = 32'h00000000 /* 0xa6c8 */;
                10675: data_o = 32'h00000000 /* 0xa6cc */;
                10676: data_o = 32'h00000000 /* 0xa6d0 */;
                10677: data_o = 32'h00000000 /* 0xa6d4 */;
                10678: data_o = 32'h00000000 /* 0xa6d8 */;
                10679: data_o = 32'h00000000 /* 0xa6dc */;
                10680: data_o = 32'h00000000 /* 0xa6e0 */;
                10681: data_o = 32'h00000000 /* 0xa6e4 */;
                10682: data_o = 32'h00000000 /* 0xa6e8 */;
                10683: data_o = 32'h00000000 /* 0xa6ec */;
                10684: data_o = 32'h00000000 /* 0xa6f0 */;
                10685: data_o = 32'h00000000 /* 0xa6f4 */;
                10686: data_o = 32'h00000000 /* 0xa6f8 */;
                10687: data_o = 32'h00000000 /* 0xa6fc */;
                10688: data_o = 32'h00000000 /* 0xa700 */;
                10689: data_o = 32'h00000000 /* 0xa704 */;
                10690: data_o = 32'h00000000 /* 0xa708 */;
                10691: data_o = 32'h00000000 /* 0xa70c */;
                10692: data_o = 32'h00000000 /* 0xa710 */;
                10693: data_o = 32'h00000000 /* 0xa714 */;
                10694: data_o = 32'h00000000 /* 0xa718 */;
                10695: data_o = 32'h00000000 /* 0xa71c */;
                10696: data_o = 32'h00000000 /* 0xa720 */;
                10697: data_o = 32'h00000000 /* 0xa724 */;
                10698: data_o = 32'h00000000 /* 0xa728 */;
                10699: data_o = 32'h00000000 /* 0xa72c */;
                10700: data_o = 32'h00000000 /* 0xa730 */;
                10701: data_o = 32'h00000000 /* 0xa734 */;
                10702: data_o = 32'h00000000 /* 0xa738 */;
                10703: data_o = 32'h00000000 /* 0xa73c */;
                10704: data_o = 32'h00000000 /* 0xa740 */;
                10705: data_o = 32'h00000000 /* 0xa744 */;
                10706: data_o = 32'h00000000 /* 0xa748 */;
                10707: data_o = 32'h00000000 /* 0xa74c */;
                10708: data_o = 32'h00000000 /* 0xa750 */;
                10709: data_o = 32'h00000000 /* 0xa754 */;
                10710: data_o = 32'h00000000 /* 0xa758 */;
                10711: data_o = 32'h00000000 /* 0xa75c */;
                10712: data_o = 32'h00000000 /* 0xa760 */;
                10713: data_o = 32'h00000000 /* 0xa764 */;
                10714: data_o = 32'h00000000 /* 0xa768 */;
                10715: data_o = 32'h00000000 /* 0xa76c */;
                10716: data_o = 32'h00000000 /* 0xa770 */;
                10717: data_o = 32'h00000000 /* 0xa774 */;
                10718: data_o = 32'h00000000 /* 0xa778 */;
                10719: data_o = 32'h00000000 /* 0xa77c */;
                10720: data_o = 32'h00000000 /* 0xa780 */;
                10721: data_o = 32'h00000000 /* 0xa784 */;
                10722: data_o = 32'h00000000 /* 0xa788 */;
                10723: data_o = 32'h00000000 /* 0xa78c */;
                10724: data_o = 32'h00000000 /* 0xa790 */;
                10725: data_o = 32'h00000000 /* 0xa794 */;
                10726: data_o = 32'h00000000 /* 0xa798 */;
                10727: data_o = 32'h00000000 /* 0xa79c */;
                10728: data_o = 32'h00000000 /* 0xa7a0 */;
                10729: data_o = 32'h00000000 /* 0xa7a4 */;
                10730: data_o = 32'h00000000 /* 0xa7a8 */;
                10731: data_o = 32'h00000000 /* 0xa7ac */;
                10732: data_o = 32'h00000000 /* 0xa7b0 */;
                10733: data_o = 32'h00000000 /* 0xa7b4 */;
                10734: data_o = 32'h00000000 /* 0xa7b8 */;
                10735: data_o = 32'h00000000 /* 0xa7bc */;
                10736: data_o = 32'h00000000 /* 0xa7c0 */;
                10737: data_o = 32'h00000000 /* 0xa7c4 */;
                10738: data_o = 32'h00000000 /* 0xa7c8 */;
                10739: data_o = 32'h00000000 /* 0xa7cc */;
                10740: data_o = 32'h00000000 /* 0xa7d0 */;
                10741: data_o = 32'h00000000 /* 0xa7d4 */;
                10742: data_o = 32'h00000000 /* 0xa7d8 */;
                10743: data_o = 32'h00000000 /* 0xa7dc */;
                10744: data_o = 32'h00000000 /* 0xa7e0 */;
                10745: data_o = 32'h00000000 /* 0xa7e4 */;
                10746: data_o = 32'h00000000 /* 0xa7e8 */;
                10747: data_o = 32'h00000000 /* 0xa7ec */;
                10748: data_o = 32'h00000000 /* 0xa7f0 */;
                10749: data_o = 32'h00000000 /* 0xa7f4 */;
                10750: data_o = 32'h00000000 /* 0xa7f8 */;
                10751: data_o = 32'h00000000 /* 0xa7fc */;
                10752: data_o = 32'h00000000 /* 0xa800 */;
                10753: data_o = 32'h00000000 /* 0xa804 */;
                10754: data_o = 32'h00000000 /* 0xa808 */;
                10755: data_o = 32'h00000000 /* 0xa80c */;
                10756: data_o = 32'h00000000 /* 0xa810 */;
                10757: data_o = 32'h00000000 /* 0xa814 */;
                10758: data_o = 32'h00000000 /* 0xa818 */;
                10759: data_o = 32'h00000000 /* 0xa81c */;
                10760: data_o = 32'h00000000 /* 0xa820 */;
                10761: data_o = 32'h00000000 /* 0xa824 */;
                10762: data_o = 32'h00000000 /* 0xa828 */;
                10763: data_o = 32'h00000000 /* 0xa82c */;
                10764: data_o = 32'h00000000 /* 0xa830 */;
                10765: data_o = 32'h00000000 /* 0xa834 */;
                10766: data_o = 32'h00000000 /* 0xa838 */;
                10767: data_o = 32'h00000000 /* 0xa83c */;
                10768: data_o = 32'h00000000 /* 0xa840 */;
                10769: data_o = 32'h00000000 /* 0xa844 */;
                10770: data_o = 32'h00000000 /* 0xa848 */;
                10771: data_o = 32'h00000000 /* 0xa84c */;
                10772: data_o = 32'h00000000 /* 0xa850 */;
                10773: data_o = 32'h00000000 /* 0xa854 */;
                10774: data_o = 32'h00000000 /* 0xa858 */;
                10775: data_o = 32'h00000000 /* 0xa85c */;
                10776: data_o = 32'h00000000 /* 0xa860 */;
                10777: data_o = 32'h00000000 /* 0xa864 */;
                10778: data_o = 32'h00000000 /* 0xa868 */;
                10779: data_o = 32'h00000000 /* 0xa86c */;
                10780: data_o = 32'h00000000 /* 0xa870 */;
                10781: data_o = 32'h00000000 /* 0xa874 */;
                10782: data_o = 32'h00000000 /* 0xa878 */;
                10783: data_o = 32'h00000000 /* 0xa87c */;
                10784: data_o = 32'h00000000 /* 0xa880 */;
                10785: data_o = 32'h00000000 /* 0xa884 */;
                10786: data_o = 32'h00000000 /* 0xa888 */;
                10787: data_o = 32'h00000000 /* 0xa88c */;
                10788: data_o = 32'h00000000 /* 0xa890 */;
                10789: data_o = 32'h00000000 /* 0xa894 */;
                10790: data_o = 32'h00000000 /* 0xa898 */;
                10791: data_o = 32'h00000000 /* 0xa89c */;
                10792: data_o = 32'h00000000 /* 0xa8a0 */;
                10793: data_o = 32'h00000000 /* 0xa8a4 */;
                10794: data_o = 32'h00000000 /* 0xa8a8 */;
                10795: data_o = 32'h00000000 /* 0xa8ac */;
                10796: data_o = 32'h00000000 /* 0xa8b0 */;
                10797: data_o = 32'h00000000 /* 0xa8b4 */;
                10798: data_o = 32'h00000000 /* 0xa8b8 */;
                10799: data_o = 32'h00000000 /* 0xa8bc */;
                10800: data_o = 32'h00000000 /* 0xa8c0 */;
                10801: data_o = 32'h00000000 /* 0xa8c4 */;
                10802: data_o = 32'h00000000 /* 0xa8c8 */;
                10803: data_o = 32'h00000000 /* 0xa8cc */;
                10804: data_o = 32'h00000000 /* 0xa8d0 */;
                10805: data_o = 32'h00000000 /* 0xa8d4 */;
                10806: data_o = 32'h00000000 /* 0xa8d8 */;
                10807: data_o = 32'h00000000 /* 0xa8dc */;
                10808: data_o = 32'h00000000 /* 0xa8e0 */;
                10809: data_o = 32'h00000000 /* 0xa8e4 */;
                10810: data_o = 32'h00000000 /* 0xa8e8 */;
                10811: data_o = 32'h00000000 /* 0xa8ec */;
                10812: data_o = 32'h00000000 /* 0xa8f0 */;
                10813: data_o = 32'h00000000 /* 0xa8f4 */;
                10814: data_o = 32'h00000000 /* 0xa8f8 */;
                10815: data_o = 32'h00000000 /* 0xa8fc */;
                10816: data_o = 32'h00000000 /* 0xa900 */;
                10817: data_o = 32'h00000000 /* 0xa904 */;
                10818: data_o = 32'h00000000 /* 0xa908 */;
                10819: data_o = 32'h00000000 /* 0xa90c */;
                10820: data_o = 32'h00000000 /* 0xa910 */;
                10821: data_o = 32'h00000000 /* 0xa914 */;
                10822: data_o = 32'h00000000 /* 0xa918 */;
                10823: data_o = 32'h00000000 /* 0xa91c */;
                10824: data_o = 32'h00000000 /* 0xa920 */;
                10825: data_o = 32'h00000000 /* 0xa924 */;
                10826: data_o = 32'h00000000 /* 0xa928 */;
                10827: data_o = 32'h00000000 /* 0xa92c */;
                10828: data_o = 32'h00000000 /* 0xa930 */;
                10829: data_o = 32'h00000000 /* 0xa934 */;
                10830: data_o = 32'h00000000 /* 0xa938 */;
                10831: data_o = 32'h00000000 /* 0xa93c */;
                10832: data_o = 32'h00000000 /* 0xa940 */;
                10833: data_o = 32'h00000000 /* 0xa944 */;
                10834: data_o = 32'h00000000 /* 0xa948 */;
                10835: data_o = 32'h00000000 /* 0xa94c */;
                10836: data_o = 32'h00000000 /* 0xa950 */;
                10837: data_o = 32'h00000000 /* 0xa954 */;
                10838: data_o = 32'h00000000 /* 0xa958 */;
                10839: data_o = 32'h00000000 /* 0xa95c */;
                10840: data_o = 32'h00000000 /* 0xa960 */;
                10841: data_o = 32'h00000000 /* 0xa964 */;
                10842: data_o = 32'h00000000 /* 0xa968 */;
                10843: data_o = 32'h00000000 /* 0xa96c */;
                10844: data_o = 32'h00000000 /* 0xa970 */;
                10845: data_o = 32'h00000000 /* 0xa974 */;
                10846: data_o = 32'h00000000 /* 0xa978 */;
                10847: data_o = 32'h00000000 /* 0xa97c */;
                10848: data_o = 32'h00000000 /* 0xa980 */;
                10849: data_o = 32'h00000000 /* 0xa984 */;
                10850: data_o = 32'h00000000 /* 0xa988 */;
                10851: data_o = 32'h00000000 /* 0xa98c */;
                10852: data_o = 32'h00000000 /* 0xa990 */;
                10853: data_o = 32'h00000000 /* 0xa994 */;
                10854: data_o = 32'h00000000 /* 0xa998 */;
                10855: data_o = 32'h00000000 /* 0xa99c */;
                10856: data_o = 32'h00000000 /* 0xa9a0 */;
                10857: data_o = 32'h00000000 /* 0xa9a4 */;
                10858: data_o = 32'h00000000 /* 0xa9a8 */;
                10859: data_o = 32'h00000000 /* 0xa9ac */;
                10860: data_o = 32'h00000000 /* 0xa9b0 */;
                10861: data_o = 32'h00000000 /* 0xa9b4 */;
                10862: data_o = 32'h00000000 /* 0xa9b8 */;
                10863: data_o = 32'h00000000 /* 0xa9bc */;
                10864: data_o = 32'h00000000 /* 0xa9c0 */;
                10865: data_o = 32'h00000000 /* 0xa9c4 */;
                10866: data_o = 32'h00000000 /* 0xa9c8 */;
                10867: data_o = 32'h00000000 /* 0xa9cc */;
                10868: data_o = 32'h00000000 /* 0xa9d0 */;
                10869: data_o = 32'h00000000 /* 0xa9d4 */;
                10870: data_o = 32'h00000000 /* 0xa9d8 */;
                10871: data_o = 32'h00000000 /* 0xa9dc */;
                10872: data_o = 32'h00000000 /* 0xa9e0 */;
                10873: data_o = 32'h00000000 /* 0xa9e4 */;
                10874: data_o = 32'h00000000 /* 0xa9e8 */;
                10875: data_o = 32'h00000000 /* 0xa9ec */;
                10876: data_o = 32'h00000000 /* 0xa9f0 */;
                10877: data_o = 32'h00000000 /* 0xa9f4 */;
                10878: data_o = 32'h00000000 /* 0xa9f8 */;
                10879: data_o = 32'h00000000 /* 0xa9fc */;
                10880: data_o = 32'h00000000 /* 0xaa00 */;
                10881: data_o = 32'h00000000 /* 0xaa04 */;
                10882: data_o = 32'h00000000 /* 0xaa08 */;
                10883: data_o = 32'h00000000 /* 0xaa0c */;
                10884: data_o = 32'h00000000 /* 0xaa10 */;
                10885: data_o = 32'h00000000 /* 0xaa14 */;
                10886: data_o = 32'h00000000 /* 0xaa18 */;
                10887: data_o = 32'h00000000 /* 0xaa1c */;
                10888: data_o = 32'h00000000 /* 0xaa20 */;
                10889: data_o = 32'h00000000 /* 0xaa24 */;
                10890: data_o = 32'h00000000 /* 0xaa28 */;
                10891: data_o = 32'h00000000 /* 0xaa2c */;
                10892: data_o = 32'h00000000 /* 0xaa30 */;
                10893: data_o = 32'h00000000 /* 0xaa34 */;
                10894: data_o = 32'h00000000 /* 0xaa38 */;
                10895: data_o = 32'h00000000 /* 0xaa3c */;
                10896: data_o = 32'h00000000 /* 0xaa40 */;
                10897: data_o = 32'h00000000 /* 0xaa44 */;
                10898: data_o = 32'h00000000 /* 0xaa48 */;
                10899: data_o = 32'h00000000 /* 0xaa4c */;
                10900: data_o = 32'h00000000 /* 0xaa50 */;
                10901: data_o = 32'h00000000 /* 0xaa54 */;
                10902: data_o = 32'h00000000 /* 0xaa58 */;
                10903: data_o = 32'h00000000 /* 0xaa5c */;
                10904: data_o = 32'h00000000 /* 0xaa60 */;
                10905: data_o = 32'h00000000 /* 0xaa64 */;
                10906: data_o = 32'h00000000 /* 0xaa68 */;
                10907: data_o = 32'h00000000 /* 0xaa6c */;
                10908: data_o = 32'h00000000 /* 0xaa70 */;
                10909: data_o = 32'h00000000 /* 0xaa74 */;
                10910: data_o = 32'h00000000 /* 0xaa78 */;
                10911: data_o = 32'h00000000 /* 0xaa7c */;
                10912: data_o = 32'h00000000 /* 0xaa80 */;
                10913: data_o = 32'h00000000 /* 0xaa84 */;
                10914: data_o = 32'h00000000 /* 0xaa88 */;
                10915: data_o = 32'h00000000 /* 0xaa8c */;
                10916: data_o = 32'h00000000 /* 0xaa90 */;
                10917: data_o = 32'h00000000 /* 0xaa94 */;
                10918: data_o = 32'h00000000 /* 0xaa98 */;
                10919: data_o = 32'h00000000 /* 0xaa9c */;
                10920: data_o = 32'h00000000 /* 0xaaa0 */;
                10921: data_o = 32'h00000000 /* 0xaaa4 */;
                10922: data_o = 32'h00000000 /* 0xaaa8 */;
                10923: data_o = 32'h00000000 /* 0xaaac */;
                10924: data_o = 32'h00000000 /* 0xaab0 */;
                10925: data_o = 32'h00000000 /* 0xaab4 */;
                10926: data_o = 32'h00000000 /* 0xaab8 */;
                10927: data_o = 32'h00000000 /* 0xaabc */;
                10928: data_o = 32'h00000000 /* 0xaac0 */;
                10929: data_o = 32'h00000000 /* 0xaac4 */;
                10930: data_o = 32'h00000000 /* 0xaac8 */;
                10931: data_o = 32'h00000000 /* 0xaacc */;
                10932: data_o = 32'h00000000 /* 0xaad0 */;
                10933: data_o = 32'h00000000 /* 0xaad4 */;
                10934: data_o = 32'h00000000 /* 0xaad8 */;
                10935: data_o = 32'h00000000 /* 0xaadc */;
                10936: data_o = 32'h00000000 /* 0xaae0 */;
                10937: data_o = 32'h00000000 /* 0xaae4 */;
                10938: data_o = 32'h00000000 /* 0xaae8 */;
                10939: data_o = 32'h00000000 /* 0xaaec */;
                10940: data_o = 32'h00000000 /* 0xaaf0 */;
                10941: data_o = 32'h00000000 /* 0xaaf4 */;
                10942: data_o = 32'h00000000 /* 0xaaf8 */;
                10943: data_o = 32'h00000000 /* 0xaafc */;
                10944: data_o = 32'h00000000 /* 0xab00 */;
                10945: data_o = 32'h00000000 /* 0xab04 */;
                10946: data_o = 32'h00000000 /* 0xab08 */;
                10947: data_o = 32'h00000000 /* 0xab0c */;
                10948: data_o = 32'h00000000 /* 0xab10 */;
                10949: data_o = 32'h00000000 /* 0xab14 */;
                10950: data_o = 32'h00000000 /* 0xab18 */;
                10951: data_o = 32'h00000000 /* 0xab1c */;
                10952: data_o = 32'h00000000 /* 0xab20 */;
                10953: data_o = 32'h00000000 /* 0xab24 */;
                10954: data_o = 32'h00000000 /* 0xab28 */;
                10955: data_o = 32'h00000000 /* 0xab2c */;
                10956: data_o = 32'h00000000 /* 0xab30 */;
                10957: data_o = 32'h00000000 /* 0xab34 */;
                10958: data_o = 32'h00000000 /* 0xab38 */;
                10959: data_o = 32'h00000000 /* 0xab3c */;
                10960: data_o = 32'h00000000 /* 0xab40 */;
                10961: data_o = 32'h00000000 /* 0xab44 */;
                10962: data_o = 32'h00000000 /* 0xab48 */;
                10963: data_o = 32'h00000000 /* 0xab4c */;
                10964: data_o = 32'h00000000 /* 0xab50 */;
                10965: data_o = 32'h00000000 /* 0xab54 */;
                10966: data_o = 32'h00000000 /* 0xab58 */;
                10967: data_o = 32'h00000000 /* 0xab5c */;
                10968: data_o = 32'h00000000 /* 0xab60 */;
                10969: data_o = 32'h00000000 /* 0xab64 */;
                10970: data_o = 32'h00000000 /* 0xab68 */;
                10971: data_o = 32'h00000000 /* 0xab6c */;
                10972: data_o = 32'h00000000 /* 0xab70 */;
                10973: data_o = 32'h00000000 /* 0xab74 */;
                10974: data_o = 32'h00000000 /* 0xab78 */;
                10975: data_o = 32'h00000000 /* 0xab7c */;
                10976: data_o = 32'h00000000 /* 0xab80 */;
                10977: data_o = 32'h00000000 /* 0xab84 */;
                10978: data_o = 32'h00000000 /* 0xab88 */;
                10979: data_o = 32'h00000000 /* 0xab8c */;
                10980: data_o = 32'h00000000 /* 0xab90 */;
                10981: data_o = 32'h00000000 /* 0xab94 */;
                10982: data_o = 32'h00000000 /* 0xab98 */;
                10983: data_o = 32'h00000000 /* 0xab9c */;
                10984: data_o = 32'h00000000 /* 0xaba0 */;
                10985: data_o = 32'h00000000 /* 0xaba4 */;
                10986: data_o = 32'h00000000 /* 0xaba8 */;
                10987: data_o = 32'h00000000 /* 0xabac */;
                10988: data_o = 32'h00000000 /* 0xabb0 */;
                10989: data_o = 32'h00000000 /* 0xabb4 */;
                10990: data_o = 32'h00000000 /* 0xabb8 */;
                10991: data_o = 32'h00000000 /* 0xabbc */;
                10992: data_o = 32'h00000000 /* 0xabc0 */;
                10993: data_o = 32'h00000000 /* 0xabc4 */;
                10994: data_o = 32'h00000000 /* 0xabc8 */;
                10995: data_o = 32'h00000000 /* 0xabcc */;
                10996: data_o = 32'h00000000 /* 0xabd0 */;
                10997: data_o = 32'h00000000 /* 0xabd4 */;
                10998: data_o = 32'h00000000 /* 0xabd8 */;
                10999: data_o = 32'h00000000 /* 0xabdc */;
                11000: data_o = 32'h00000000 /* 0xabe0 */;
                11001: data_o = 32'h00000000 /* 0xabe4 */;
                11002: data_o = 32'h00000000 /* 0xabe8 */;
                11003: data_o = 32'h00000000 /* 0xabec */;
                11004: data_o = 32'h00000000 /* 0xabf0 */;
                11005: data_o = 32'h00000000 /* 0xabf4 */;
                11006: data_o = 32'h00000000 /* 0xabf8 */;
                11007: data_o = 32'h00000000 /* 0xabfc */;
                11008: data_o = 32'h00000000 /* 0xac00 */;
                11009: data_o = 32'h00000000 /* 0xac04 */;
                11010: data_o = 32'h00000000 /* 0xac08 */;
                11011: data_o = 32'h00000000 /* 0xac0c */;
                11012: data_o = 32'h00000000 /* 0xac10 */;
                11013: data_o = 32'h00000000 /* 0xac14 */;
                11014: data_o = 32'h00000000 /* 0xac18 */;
                11015: data_o = 32'h00000000 /* 0xac1c */;
                11016: data_o = 32'h00000000 /* 0xac20 */;
                11017: data_o = 32'h00000000 /* 0xac24 */;
                11018: data_o = 32'h00000000 /* 0xac28 */;
                11019: data_o = 32'h00000000 /* 0xac2c */;
                11020: data_o = 32'h00000000 /* 0xac30 */;
                11021: data_o = 32'h00000000 /* 0xac34 */;
                11022: data_o = 32'h00000000 /* 0xac38 */;
                11023: data_o = 32'h00000000 /* 0xac3c */;
                11024: data_o = 32'h00000000 /* 0xac40 */;
                11025: data_o = 32'h00000000 /* 0xac44 */;
                11026: data_o = 32'h00000000 /* 0xac48 */;
                11027: data_o = 32'h00000000 /* 0xac4c */;
                11028: data_o = 32'h00000000 /* 0xac50 */;
                11029: data_o = 32'h00000000 /* 0xac54 */;
                11030: data_o = 32'h00000000 /* 0xac58 */;
                11031: data_o = 32'h00000000 /* 0xac5c */;
                11032: data_o = 32'h00000000 /* 0xac60 */;
                11033: data_o = 32'h00000000 /* 0xac64 */;
                11034: data_o = 32'h00000000 /* 0xac68 */;
                11035: data_o = 32'h00000000 /* 0xac6c */;
                11036: data_o = 32'h00000000 /* 0xac70 */;
                11037: data_o = 32'h00000000 /* 0xac74 */;
                11038: data_o = 32'h00000000 /* 0xac78 */;
                11039: data_o = 32'h00000000 /* 0xac7c */;
                11040: data_o = 32'h00000000 /* 0xac80 */;
                11041: data_o = 32'h00000000 /* 0xac84 */;
                11042: data_o = 32'h00000000 /* 0xac88 */;
                11043: data_o = 32'h00000000 /* 0xac8c */;
                11044: data_o = 32'h00000000 /* 0xac90 */;
                11045: data_o = 32'h00000000 /* 0xac94 */;
                11046: data_o = 32'h00000000 /* 0xac98 */;
                11047: data_o = 32'h00000000 /* 0xac9c */;
                11048: data_o = 32'h00000000 /* 0xaca0 */;
                11049: data_o = 32'h00000000 /* 0xaca4 */;
                11050: data_o = 32'h00000000 /* 0xaca8 */;
                11051: data_o = 32'h00000000 /* 0xacac */;
                11052: data_o = 32'h00000000 /* 0xacb0 */;
                11053: data_o = 32'h00000000 /* 0xacb4 */;
                11054: data_o = 32'h00000000 /* 0xacb8 */;
                11055: data_o = 32'h00000000 /* 0xacbc */;
                11056: data_o = 32'h00000000 /* 0xacc0 */;
                11057: data_o = 32'h00000000 /* 0xacc4 */;
                11058: data_o = 32'h00000000 /* 0xacc8 */;
                11059: data_o = 32'h00000000 /* 0xaccc */;
                11060: data_o = 32'h00000000 /* 0xacd0 */;
                11061: data_o = 32'h00000000 /* 0xacd4 */;
                11062: data_o = 32'h00000000 /* 0xacd8 */;
                11063: data_o = 32'h00000000 /* 0xacdc */;
                11064: data_o = 32'h00000000 /* 0xace0 */;
                11065: data_o = 32'h00000000 /* 0xace4 */;
                11066: data_o = 32'h00000000 /* 0xace8 */;
                11067: data_o = 32'h00000000 /* 0xacec */;
                11068: data_o = 32'h00000000 /* 0xacf0 */;
                11069: data_o = 32'h00000000 /* 0xacf4 */;
                11070: data_o = 32'h00000000 /* 0xacf8 */;
                11071: data_o = 32'h00000000 /* 0xacfc */;
                11072: data_o = 32'h00000000 /* 0xad00 */;
                11073: data_o = 32'h00000000 /* 0xad04 */;
                11074: data_o = 32'h00000000 /* 0xad08 */;
                11075: data_o = 32'h00000000 /* 0xad0c */;
                11076: data_o = 32'h00000000 /* 0xad10 */;
                11077: data_o = 32'h00000000 /* 0xad14 */;
                11078: data_o = 32'h00000000 /* 0xad18 */;
                11079: data_o = 32'h00000000 /* 0xad1c */;
                11080: data_o = 32'h00000000 /* 0xad20 */;
                11081: data_o = 32'h00000000 /* 0xad24 */;
                11082: data_o = 32'h00000000 /* 0xad28 */;
                11083: data_o = 32'h00000000 /* 0xad2c */;
                11084: data_o = 32'h00000000 /* 0xad30 */;
                11085: data_o = 32'h00000000 /* 0xad34 */;
                11086: data_o = 32'h00000000 /* 0xad38 */;
                11087: data_o = 32'h00000000 /* 0xad3c */;
                11088: data_o = 32'h00000000 /* 0xad40 */;
                11089: data_o = 32'h00000000 /* 0xad44 */;
                11090: data_o = 32'h00000000 /* 0xad48 */;
                11091: data_o = 32'h00000000 /* 0xad4c */;
                11092: data_o = 32'h00000000 /* 0xad50 */;
                11093: data_o = 32'h00000000 /* 0xad54 */;
                11094: data_o = 32'h00000000 /* 0xad58 */;
                11095: data_o = 32'h00000000 /* 0xad5c */;
                11096: data_o = 32'h00000000 /* 0xad60 */;
                11097: data_o = 32'h00000000 /* 0xad64 */;
                11098: data_o = 32'h00000000 /* 0xad68 */;
                11099: data_o = 32'h00000000 /* 0xad6c */;
                11100: data_o = 32'h00000000 /* 0xad70 */;
                11101: data_o = 32'h00000000 /* 0xad74 */;
                11102: data_o = 32'h00000000 /* 0xad78 */;
                11103: data_o = 32'h00000000 /* 0xad7c */;
                11104: data_o = 32'h00000000 /* 0xad80 */;
                11105: data_o = 32'h00000000 /* 0xad84 */;
                11106: data_o = 32'h00000000 /* 0xad88 */;
                11107: data_o = 32'h00000000 /* 0xad8c */;
                11108: data_o = 32'h00000000 /* 0xad90 */;
                11109: data_o = 32'h00000000 /* 0xad94 */;
                11110: data_o = 32'h00000000 /* 0xad98 */;
                11111: data_o = 32'h00000000 /* 0xad9c */;
                11112: data_o = 32'h00000000 /* 0xada0 */;
                11113: data_o = 32'h00000000 /* 0xada4 */;
                11114: data_o = 32'h00000000 /* 0xada8 */;
                11115: data_o = 32'h00000000 /* 0xadac */;
                11116: data_o = 32'h00000000 /* 0xadb0 */;
                11117: data_o = 32'h00000000 /* 0xadb4 */;
                11118: data_o = 32'h00000000 /* 0xadb8 */;
                11119: data_o = 32'h00000000 /* 0xadbc */;
                11120: data_o = 32'h00000000 /* 0xadc0 */;
                11121: data_o = 32'h00000000 /* 0xadc4 */;
                11122: data_o = 32'h00000000 /* 0xadc8 */;
                11123: data_o = 32'h00000000 /* 0xadcc */;
                11124: data_o = 32'h00000000 /* 0xadd0 */;
                11125: data_o = 32'h00000000 /* 0xadd4 */;
                11126: data_o = 32'h00000000 /* 0xadd8 */;
                11127: data_o = 32'h00000000 /* 0xaddc */;
                11128: data_o = 32'h00000000 /* 0xade0 */;
                11129: data_o = 32'h00000000 /* 0xade4 */;
                11130: data_o = 32'h00000000 /* 0xade8 */;
                11131: data_o = 32'h00000000 /* 0xadec */;
                11132: data_o = 32'h00000000 /* 0xadf0 */;
                11133: data_o = 32'h00000000 /* 0xadf4 */;
                11134: data_o = 32'h00000000 /* 0xadf8 */;
                11135: data_o = 32'h00000000 /* 0xadfc */;
                11136: data_o = 32'h00000000 /* 0xae00 */;
                11137: data_o = 32'h00000000 /* 0xae04 */;
                11138: data_o = 32'h00000000 /* 0xae08 */;
                11139: data_o = 32'h00000000 /* 0xae0c */;
                11140: data_o = 32'h00000000 /* 0xae10 */;
                11141: data_o = 32'h00000000 /* 0xae14 */;
                11142: data_o = 32'h00000000 /* 0xae18 */;
                11143: data_o = 32'h00000000 /* 0xae1c */;
                11144: data_o = 32'h00000000 /* 0xae20 */;
                11145: data_o = 32'h00000000 /* 0xae24 */;
                11146: data_o = 32'h00000000 /* 0xae28 */;
                11147: data_o = 32'h00000000 /* 0xae2c */;
                11148: data_o = 32'h00000000 /* 0xae30 */;
                11149: data_o = 32'h00000000 /* 0xae34 */;
                11150: data_o = 32'h00000000 /* 0xae38 */;
                11151: data_o = 32'h00000000 /* 0xae3c */;
                11152: data_o = 32'h00000000 /* 0xae40 */;
                11153: data_o = 32'h00000000 /* 0xae44 */;
                11154: data_o = 32'h00000000 /* 0xae48 */;
                11155: data_o = 32'h00000000 /* 0xae4c */;
                11156: data_o = 32'h00000000 /* 0xae50 */;
                11157: data_o = 32'h00000000 /* 0xae54 */;
                11158: data_o = 32'h00000000 /* 0xae58 */;
                11159: data_o = 32'h00000000 /* 0xae5c */;
                11160: data_o = 32'h00000000 /* 0xae60 */;
                11161: data_o = 32'h00000000 /* 0xae64 */;
                11162: data_o = 32'h00000000 /* 0xae68 */;
                11163: data_o = 32'h00000000 /* 0xae6c */;
                11164: data_o = 32'h00000000 /* 0xae70 */;
                11165: data_o = 32'h00000000 /* 0xae74 */;
                11166: data_o = 32'h00000000 /* 0xae78 */;
                11167: data_o = 32'h00000000 /* 0xae7c */;
                11168: data_o = 32'h00000000 /* 0xae80 */;
                11169: data_o = 32'h00000000 /* 0xae84 */;
                11170: data_o = 32'h00000000 /* 0xae88 */;
                11171: data_o = 32'h00000000 /* 0xae8c */;
                11172: data_o = 32'h00000000 /* 0xae90 */;
                11173: data_o = 32'h00000000 /* 0xae94 */;
                11174: data_o = 32'h00000000 /* 0xae98 */;
                11175: data_o = 32'h00000000 /* 0xae9c */;
                11176: data_o = 32'h00000000 /* 0xaea0 */;
                11177: data_o = 32'h00000000 /* 0xaea4 */;
                11178: data_o = 32'h00000000 /* 0xaea8 */;
                11179: data_o = 32'h00000000 /* 0xaeac */;
                11180: data_o = 32'h00000000 /* 0xaeb0 */;
                11181: data_o = 32'h00000000 /* 0xaeb4 */;
                11182: data_o = 32'h00000000 /* 0xaeb8 */;
                11183: data_o = 32'h00000000 /* 0xaebc */;
                11184: data_o = 32'h00000000 /* 0xaec0 */;
                11185: data_o = 32'h00000000 /* 0xaec4 */;
                11186: data_o = 32'h00000000 /* 0xaec8 */;
                11187: data_o = 32'h00000000 /* 0xaecc */;
                11188: data_o = 32'h00000000 /* 0xaed0 */;
                11189: data_o = 32'h00000000 /* 0xaed4 */;
                11190: data_o = 32'h00000000 /* 0xaed8 */;
                11191: data_o = 32'h00000000 /* 0xaedc */;
                11192: data_o = 32'h00000000 /* 0xaee0 */;
                11193: data_o = 32'h00000000 /* 0xaee4 */;
                11194: data_o = 32'h00000000 /* 0xaee8 */;
                11195: data_o = 32'h00000000 /* 0xaeec */;
                11196: data_o = 32'h00000000 /* 0xaef0 */;
                11197: data_o = 32'h00000000 /* 0xaef4 */;
                11198: data_o = 32'h00000000 /* 0xaef8 */;
                11199: data_o = 32'h00000000 /* 0xaefc */;
                11200: data_o = 32'h00000000 /* 0xaf00 */;
                11201: data_o = 32'h00000000 /* 0xaf04 */;
                11202: data_o = 32'h00000000 /* 0xaf08 */;
                11203: data_o = 32'h00000000 /* 0xaf0c */;
                11204: data_o = 32'h00000000 /* 0xaf10 */;
                11205: data_o = 32'h00000000 /* 0xaf14 */;
                11206: data_o = 32'h00000000 /* 0xaf18 */;
                11207: data_o = 32'h00000000 /* 0xaf1c */;
                11208: data_o = 32'h00000000 /* 0xaf20 */;
                11209: data_o = 32'h00000000 /* 0xaf24 */;
                11210: data_o = 32'h00000000 /* 0xaf28 */;
                11211: data_o = 32'h00000000 /* 0xaf2c */;
                11212: data_o = 32'h00000000 /* 0xaf30 */;
                11213: data_o = 32'h00000000 /* 0xaf34 */;
                11214: data_o = 32'h00000000 /* 0xaf38 */;
                11215: data_o = 32'h00000000 /* 0xaf3c */;
                11216: data_o = 32'h00000000 /* 0xaf40 */;
                11217: data_o = 32'h00000000 /* 0xaf44 */;
                11218: data_o = 32'h00000000 /* 0xaf48 */;
                11219: data_o = 32'h00000000 /* 0xaf4c */;
                11220: data_o = 32'h00000000 /* 0xaf50 */;
                11221: data_o = 32'h00000000 /* 0xaf54 */;
                11222: data_o = 32'h00000000 /* 0xaf58 */;
                11223: data_o = 32'h00000000 /* 0xaf5c */;
                11224: data_o = 32'h00000000 /* 0xaf60 */;
                11225: data_o = 32'h00000000 /* 0xaf64 */;
                11226: data_o = 32'h00000000 /* 0xaf68 */;
                11227: data_o = 32'h00000000 /* 0xaf6c */;
                11228: data_o = 32'h00000000 /* 0xaf70 */;
                11229: data_o = 32'h00000000 /* 0xaf74 */;
                11230: data_o = 32'h00000000 /* 0xaf78 */;
                11231: data_o = 32'h00000000 /* 0xaf7c */;
                11232: data_o = 32'h00000000 /* 0xaf80 */;
                11233: data_o = 32'h00000000 /* 0xaf84 */;
                11234: data_o = 32'h00000000 /* 0xaf88 */;
                11235: data_o = 32'h00000000 /* 0xaf8c */;
                11236: data_o = 32'h00000000 /* 0xaf90 */;
                11237: data_o = 32'h00000000 /* 0xaf94 */;
                11238: data_o = 32'h00000000 /* 0xaf98 */;
                11239: data_o = 32'h00000000 /* 0xaf9c */;
                11240: data_o = 32'h00000000 /* 0xafa0 */;
                11241: data_o = 32'h00000000 /* 0xafa4 */;
                11242: data_o = 32'h00000000 /* 0xafa8 */;
                11243: data_o = 32'h00000000 /* 0xafac */;
                11244: data_o = 32'h00000000 /* 0xafb0 */;
                11245: data_o = 32'h00000000 /* 0xafb4 */;
                11246: data_o = 32'h00000000 /* 0xafb8 */;
                11247: data_o = 32'h00000000 /* 0xafbc */;
                11248: data_o = 32'h00000000 /* 0xafc0 */;
                11249: data_o = 32'h00000000 /* 0xafc4 */;
                11250: data_o = 32'h00000000 /* 0xafc8 */;
                11251: data_o = 32'h00000000 /* 0xafcc */;
                11252: data_o = 32'h00000000 /* 0xafd0 */;
                11253: data_o = 32'h00000000 /* 0xafd4 */;
                11254: data_o = 32'h00000000 /* 0xafd8 */;
                11255: data_o = 32'h00000000 /* 0xafdc */;
                11256: data_o = 32'h00000000 /* 0xafe0 */;
                11257: data_o = 32'h00000000 /* 0xafe4 */;
                11258: data_o = 32'h00000000 /* 0xafe8 */;
                11259: data_o = 32'h00000000 /* 0xafec */;
                11260: data_o = 32'h00000000 /* 0xaff0 */;
                11261: data_o = 32'h00000000 /* 0xaff4 */;
                11262: data_o = 32'h00000000 /* 0xaff8 */;
                11263: data_o = 32'h00000000 /* 0xaffc */;
                11264: data_o = 32'h00000000 /* 0xb000 */;
                11265: data_o = 32'h00000000 /* 0xb004 */;
                11266: data_o = 32'h00000000 /* 0xb008 */;
                11267: data_o = 32'h00000000 /* 0xb00c */;
                11268: data_o = 32'h00000000 /* 0xb010 */;
                11269: data_o = 32'h00000000 /* 0xb014 */;
                11270: data_o = 32'h00000000 /* 0xb018 */;
                11271: data_o = 32'h00000000 /* 0xb01c */;
                11272: data_o = 32'h00000000 /* 0xb020 */;
                11273: data_o = 32'h00000000 /* 0xb024 */;
                11274: data_o = 32'h00000000 /* 0xb028 */;
                11275: data_o = 32'h00000000 /* 0xb02c */;
                11276: data_o = 32'h00000000 /* 0xb030 */;
                11277: data_o = 32'h00000000 /* 0xb034 */;
                11278: data_o = 32'h00000000 /* 0xb038 */;
                11279: data_o = 32'h00000000 /* 0xb03c */;
                11280: data_o = 32'h00000000 /* 0xb040 */;
                11281: data_o = 32'h00000000 /* 0xb044 */;
                11282: data_o = 32'h00000000 /* 0xb048 */;
                11283: data_o = 32'h00000000 /* 0xb04c */;
                11284: data_o = 32'h00000000 /* 0xb050 */;
                11285: data_o = 32'h00000000 /* 0xb054 */;
                11286: data_o = 32'h00000000 /* 0xb058 */;
                11287: data_o = 32'h00000000 /* 0xb05c */;
                11288: data_o = 32'h00000000 /* 0xb060 */;
                11289: data_o = 32'h00000000 /* 0xb064 */;
                11290: data_o = 32'h00000000 /* 0xb068 */;
                11291: data_o = 32'h00000000 /* 0xb06c */;
                11292: data_o = 32'h00000000 /* 0xb070 */;
                11293: data_o = 32'h00000000 /* 0xb074 */;
                11294: data_o = 32'h00000000 /* 0xb078 */;
                11295: data_o = 32'h00000000 /* 0xb07c */;
                11296: data_o = 32'h00000000 /* 0xb080 */;
                11297: data_o = 32'h00000000 /* 0xb084 */;
                11298: data_o = 32'h00000000 /* 0xb088 */;
                11299: data_o = 32'h00000000 /* 0xb08c */;
                11300: data_o = 32'h00000000 /* 0xb090 */;
                11301: data_o = 32'h00000000 /* 0xb094 */;
                11302: data_o = 32'h00000000 /* 0xb098 */;
                11303: data_o = 32'h00000000 /* 0xb09c */;
                11304: data_o = 32'h00000000 /* 0xb0a0 */;
                11305: data_o = 32'h00000000 /* 0xb0a4 */;
                11306: data_o = 32'h00000000 /* 0xb0a8 */;
                11307: data_o = 32'h00000000 /* 0xb0ac */;
                11308: data_o = 32'h00000000 /* 0xb0b0 */;
                11309: data_o = 32'h00000000 /* 0xb0b4 */;
                11310: data_o = 32'h00000000 /* 0xb0b8 */;
                11311: data_o = 32'h00000000 /* 0xb0bc */;
                11312: data_o = 32'h00000000 /* 0xb0c0 */;
                11313: data_o = 32'h00000000 /* 0xb0c4 */;
                11314: data_o = 32'h00000000 /* 0xb0c8 */;
                11315: data_o = 32'h00000000 /* 0xb0cc */;
                11316: data_o = 32'h00000000 /* 0xb0d0 */;
                11317: data_o = 32'h00000000 /* 0xb0d4 */;
                11318: data_o = 32'h00000000 /* 0xb0d8 */;
                11319: data_o = 32'h00000000 /* 0xb0dc */;
                11320: data_o = 32'h00000000 /* 0xb0e0 */;
                11321: data_o = 32'h00000000 /* 0xb0e4 */;
                11322: data_o = 32'h00000000 /* 0xb0e8 */;
                11323: data_o = 32'h00000000 /* 0xb0ec */;
                11324: data_o = 32'h00000000 /* 0xb0f0 */;
                11325: data_o = 32'h00000000 /* 0xb0f4 */;
                11326: data_o = 32'h00000000 /* 0xb0f8 */;
                11327: data_o = 32'h00000000 /* 0xb0fc */;
                11328: data_o = 32'h00000000 /* 0xb100 */;
                11329: data_o = 32'h00000000 /* 0xb104 */;
                11330: data_o = 32'h00000000 /* 0xb108 */;
                11331: data_o = 32'h00000000 /* 0xb10c */;
                11332: data_o = 32'h00000000 /* 0xb110 */;
                11333: data_o = 32'h00000000 /* 0xb114 */;
                11334: data_o = 32'h00000000 /* 0xb118 */;
                11335: data_o = 32'h00000000 /* 0xb11c */;
                11336: data_o = 32'h00000000 /* 0xb120 */;
                11337: data_o = 32'h00000000 /* 0xb124 */;
                11338: data_o = 32'h00000000 /* 0xb128 */;
                11339: data_o = 32'h00000000 /* 0xb12c */;
                11340: data_o = 32'h00000000 /* 0xb130 */;
                11341: data_o = 32'h00000000 /* 0xb134 */;
                11342: data_o = 32'h00000000 /* 0xb138 */;
                11343: data_o = 32'h00000000 /* 0xb13c */;
                11344: data_o = 32'h00000000 /* 0xb140 */;
                11345: data_o = 32'h00000000 /* 0xb144 */;
                11346: data_o = 32'h00000000 /* 0xb148 */;
                11347: data_o = 32'h00000000 /* 0xb14c */;
                11348: data_o = 32'h00000000 /* 0xb150 */;
                11349: data_o = 32'h00000000 /* 0xb154 */;
                11350: data_o = 32'h00000000 /* 0xb158 */;
                11351: data_o = 32'h00000000 /* 0xb15c */;
                11352: data_o = 32'h00000000 /* 0xb160 */;
                11353: data_o = 32'h00000000 /* 0xb164 */;
                11354: data_o = 32'h00000000 /* 0xb168 */;
                11355: data_o = 32'h00000000 /* 0xb16c */;
                11356: data_o = 32'h00000000 /* 0xb170 */;
                11357: data_o = 32'h00000000 /* 0xb174 */;
                11358: data_o = 32'h00000000 /* 0xb178 */;
                11359: data_o = 32'h00000000 /* 0xb17c */;
                11360: data_o = 32'h00000000 /* 0xb180 */;
                11361: data_o = 32'h00000000 /* 0xb184 */;
                11362: data_o = 32'h00000000 /* 0xb188 */;
                11363: data_o = 32'h00000000 /* 0xb18c */;
                11364: data_o = 32'h00000000 /* 0xb190 */;
                11365: data_o = 32'h00000000 /* 0xb194 */;
                11366: data_o = 32'h00000000 /* 0xb198 */;
                11367: data_o = 32'h00000000 /* 0xb19c */;
                11368: data_o = 32'h00000000 /* 0xb1a0 */;
                11369: data_o = 32'h00000000 /* 0xb1a4 */;
                11370: data_o = 32'h00000000 /* 0xb1a8 */;
                11371: data_o = 32'h00000000 /* 0xb1ac */;
                11372: data_o = 32'h00000000 /* 0xb1b0 */;
                11373: data_o = 32'h00000000 /* 0xb1b4 */;
                11374: data_o = 32'h00000000 /* 0xb1b8 */;
                11375: data_o = 32'h00000000 /* 0xb1bc */;
                11376: data_o = 32'h00000000 /* 0xb1c0 */;
                11377: data_o = 32'h00000000 /* 0xb1c4 */;
                11378: data_o = 32'h00000000 /* 0xb1c8 */;
                11379: data_o = 32'h00000000 /* 0xb1cc */;
                11380: data_o = 32'h00000000 /* 0xb1d0 */;
                11381: data_o = 32'h00000000 /* 0xb1d4 */;
                11382: data_o = 32'h00000000 /* 0xb1d8 */;
                11383: data_o = 32'h00000000 /* 0xb1dc */;
                11384: data_o = 32'h00000000 /* 0xb1e0 */;
                11385: data_o = 32'h00000000 /* 0xb1e4 */;
                11386: data_o = 32'h00000000 /* 0xb1e8 */;
                11387: data_o = 32'h00000000 /* 0xb1ec */;
                11388: data_o = 32'h00000000 /* 0xb1f0 */;
                11389: data_o = 32'h00000000 /* 0xb1f4 */;
                11390: data_o = 32'h00000000 /* 0xb1f8 */;
                11391: data_o = 32'h00000000 /* 0xb1fc */;
                11392: data_o = 32'h00000000 /* 0xb200 */;
                11393: data_o = 32'h00000000 /* 0xb204 */;
                11394: data_o = 32'h00000000 /* 0xb208 */;
                11395: data_o = 32'h00000000 /* 0xb20c */;
                11396: data_o = 32'h00000000 /* 0xb210 */;
                11397: data_o = 32'h00000000 /* 0xb214 */;
                11398: data_o = 32'h00000000 /* 0xb218 */;
                11399: data_o = 32'h00000000 /* 0xb21c */;
                11400: data_o = 32'h00000000 /* 0xb220 */;
                11401: data_o = 32'h00000000 /* 0xb224 */;
                11402: data_o = 32'h00000000 /* 0xb228 */;
                11403: data_o = 32'h00000000 /* 0xb22c */;
                11404: data_o = 32'h00000000 /* 0xb230 */;
                11405: data_o = 32'h00000000 /* 0xb234 */;
                11406: data_o = 32'h00000000 /* 0xb238 */;
                11407: data_o = 32'h00000000 /* 0xb23c */;
                11408: data_o = 32'h00000000 /* 0xb240 */;
                11409: data_o = 32'h00000000 /* 0xb244 */;
                11410: data_o = 32'h00000000 /* 0xb248 */;
                11411: data_o = 32'h00000000 /* 0xb24c */;
                11412: data_o = 32'h00000000 /* 0xb250 */;
                11413: data_o = 32'h00000000 /* 0xb254 */;
                11414: data_o = 32'h00000000 /* 0xb258 */;
                11415: data_o = 32'h00000000 /* 0xb25c */;
                11416: data_o = 32'h00000000 /* 0xb260 */;
                11417: data_o = 32'h00000000 /* 0xb264 */;
                11418: data_o = 32'h00000000 /* 0xb268 */;
                11419: data_o = 32'h00000000 /* 0xb26c */;
                11420: data_o = 32'h00000000 /* 0xb270 */;
                11421: data_o = 32'h00000000 /* 0xb274 */;
                11422: data_o = 32'h00000000 /* 0xb278 */;
                11423: data_o = 32'h00000000 /* 0xb27c */;
                11424: data_o = 32'h00000000 /* 0xb280 */;
                11425: data_o = 32'h00000000 /* 0xb284 */;
                11426: data_o = 32'h00000000 /* 0xb288 */;
                11427: data_o = 32'h00000000 /* 0xb28c */;
                11428: data_o = 32'h00000000 /* 0xb290 */;
                11429: data_o = 32'h00000000 /* 0xb294 */;
                11430: data_o = 32'h00000000 /* 0xb298 */;
                11431: data_o = 32'h00000000 /* 0xb29c */;
                11432: data_o = 32'h00000000 /* 0xb2a0 */;
                11433: data_o = 32'h00000000 /* 0xb2a4 */;
                11434: data_o = 32'h00000000 /* 0xb2a8 */;
                11435: data_o = 32'h00000000 /* 0xb2ac */;
                11436: data_o = 32'h00000000 /* 0xb2b0 */;
                11437: data_o = 32'h00000000 /* 0xb2b4 */;
                11438: data_o = 32'h00000000 /* 0xb2b8 */;
                11439: data_o = 32'h00000000 /* 0xb2bc */;
                11440: data_o = 32'h00000000 /* 0xb2c0 */;
                11441: data_o = 32'h00000000 /* 0xb2c4 */;
                11442: data_o = 32'h00000000 /* 0xb2c8 */;
                11443: data_o = 32'h00000000 /* 0xb2cc */;
                11444: data_o = 32'h00000000 /* 0xb2d0 */;
                11445: data_o = 32'h00000000 /* 0xb2d4 */;
                11446: data_o = 32'h00000000 /* 0xb2d8 */;
                11447: data_o = 32'h00000000 /* 0xb2dc */;
                11448: data_o = 32'h00000000 /* 0xb2e0 */;
                11449: data_o = 32'h00000000 /* 0xb2e4 */;
                11450: data_o = 32'h00000000 /* 0xb2e8 */;
                11451: data_o = 32'h00000000 /* 0xb2ec */;
                11452: data_o = 32'h00000000 /* 0xb2f0 */;
                11453: data_o = 32'h00000000 /* 0xb2f4 */;
                11454: data_o = 32'h00000000 /* 0xb2f8 */;
                11455: data_o = 32'h00000000 /* 0xb2fc */;
                11456: data_o = 32'h00000000 /* 0xb300 */;
                11457: data_o = 32'h00000000 /* 0xb304 */;
                11458: data_o = 32'h00000000 /* 0xb308 */;
                11459: data_o = 32'h00000000 /* 0xb30c */;
                11460: data_o = 32'h00000000 /* 0xb310 */;
                11461: data_o = 32'h00000000 /* 0xb314 */;
                11462: data_o = 32'h00000000 /* 0xb318 */;
                11463: data_o = 32'h00000000 /* 0xb31c */;
                11464: data_o = 32'h00000000 /* 0xb320 */;
                11465: data_o = 32'h00000000 /* 0xb324 */;
                11466: data_o = 32'h00000000 /* 0xb328 */;
                11467: data_o = 32'h00000000 /* 0xb32c */;
                11468: data_o = 32'h00000000 /* 0xb330 */;
                11469: data_o = 32'h00000000 /* 0xb334 */;
                11470: data_o = 32'h00000000 /* 0xb338 */;
                11471: data_o = 32'h00000000 /* 0xb33c */;
                11472: data_o = 32'h00000000 /* 0xb340 */;
                11473: data_o = 32'h00000000 /* 0xb344 */;
                11474: data_o = 32'h00000000 /* 0xb348 */;
                11475: data_o = 32'h00000000 /* 0xb34c */;
                11476: data_o = 32'h00000000 /* 0xb350 */;
                11477: data_o = 32'h00000000 /* 0xb354 */;
                11478: data_o = 32'h00000000 /* 0xb358 */;
                11479: data_o = 32'h00000000 /* 0xb35c */;
                11480: data_o = 32'h00000000 /* 0xb360 */;
                11481: data_o = 32'h00000000 /* 0xb364 */;
                11482: data_o = 32'h00000000 /* 0xb368 */;
                11483: data_o = 32'h00000000 /* 0xb36c */;
                11484: data_o = 32'h00000000 /* 0xb370 */;
                11485: data_o = 32'h00000000 /* 0xb374 */;
                11486: data_o = 32'h00000000 /* 0xb378 */;
                11487: data_o = 32'h00000000 /* 0xb37c */;
                11488: data_o = 32'h00000000 /* 0xb380 */;
                11489: data_o = 32'h00000000 /* 0xb384 */;
                11490: data_o = 32'h00000000 /* 0xb388 */;
                11491: data_o = 32'h00000000 /* 0xb38c */;
                11492: data_o = 32'h00000000 /* 0xb390 */;
                11493: data_o = 32'h00000000 /* 0xb394 */;
                11494: data_o = 32'h00000000 /* 0xb398 */;
                11495: data_o = 32'h00000000 /* 0xb39c */;
                11496: data_o = 32'h00000000 /* 0xb3a0 */;
                11497: data_o = 32'h00000000 /* 0xb3a4 */;
                11498: data_o = 32'h00000000 /* 0xb3a8 */;
                11499: data_o = 32'h00000000 /* 0xb3ac */;
                11500: data_o = 32'h00000000 /* 0xb3b0 */;
                11501: data_o = 32'h00000000 /* 0xb3b4 */;
                11502: data_o = 32'h00000000 /* 0xb3b8 */;
                11503: data_o = 32'h00000000 /* 0xb3bc */;
                11504: data_o = 32'h00000000 /* 0xb3c0 */;
                11505: data_o = 32'h00000000 /* 0xb3c4 */;
                11506: data_o = 32'h00000000 /* 0xb3c8 */;
                11507: data_o = 32'h00000000 /* 0xb3cc */;
                11508: data_o = 32'h00000000 /* 0xb3d0 */;
                11509: data_o = 32'h00000000 /* 0xb3d4 */;
                11510: data_o = 32'h00000000 /* 0xb3d8 */;
                11511: data_o = 32'h00000000 /* 0xb3dc */;
                11512: data_o = 32'h00000000 /* 0xb3e0 */;
                11513: data_o = 32'h00000000 /* 0xb3e4 */;
                11514: data_o = 32'h00000000 /* 0xb3e8 */;
                11515: data_o = 32'h00000000 /* 0xb3ec */;
                11516: data_o = 32'h00000000 /* 0xb3f0 */;
                11517: data_o = 32'h00000000 /* 0xb3f4 */;
                11518: data_o = 32'h00000000 /* 0xb3f8 */;
                11519: data_o = 32'h00000000 /* 0xb3fc */;
                11520: data_o = 32'h00000000 /* 0xb400 */;
                11521: data_o = 32'h00000000 /* 0xb404 */;
                11522: data_o = 32'h00000000 /* 0xb408 */;
                11523: data_o = 32'h00000000 /* 0xb40c */;
                11524: data_o = 32'h00000000 /* 0xb410 */;
                11525: data_o = 32'h00000000 /* 0xb414 */;
                11526: data_o = 32'h00000000 /* 0xb418 */;
                11527: data_o = 32'h00000000 /* 0xb41c */;
                11528: data_o = 32'h00000000 /* 0xb420 */;
                11529: data_o = 32'h00000000 /* 0xb424 */;
                11530: data_o = 32'h00000000 /* 0xb428 */;
                11531: data_o = 32'h00000000 /* 0xb42c */;
                11532: data_o = 32'h00000000 /* 0xb430 */;
                11533: data_o = 32'h00000000 /* 0xb434 */;
                11534: data_o = 32'h00000000 /* 0xb438 */;
                11535: data_o = 32'h00000000 /* 0xb43c */;
                11536: data_o = 32'h00000000 /* 0xb440 */;
                11537: data_o = 32'h00000000 /* 0xb444 */;
                11538: data_o = 32'h00000000 /* 0xb448 */;
                11539: data_o = 32'h00000000 /* 0xb44c */;
                11540: data_o = 32'h00000000 /* 0xb450 */;
                11541: data_o = 32'h00000000 /* 0xb454 */;
                11542: data_o = 32'h00000000 /* 0xb458 */;
                11543: data_o = 32'h00000000 /* 0xb45c */;
                11544: data_o = 32'h00000000 /* 0xb460 */;
                11545: data_o = 32'h00000000 /* 0xb464 */;
                11546: data_o = 32'h00000000 /* 0xb468 */;
                11547: data_o = 32'h00000000 /* 0xb46c */;
                11548: data_o = 32'h00000000 /* 0xb470 */;
                11549: data_o = 32'h00000000 /* 0xb474 */;
                11550: data_o = 32'h00000000 /* 0xb478 */;
                11551: data_o = 32'h00000000 /* 0xb47c */;
                11552: data_o = 32'h00000000 /* 0xb480 */;
                11553: data_o = 32'h00000000 /* 0xb484 */;
                11554: data_o = 32'h00000000 /* 0xb488 */;
                11555: data_o = 32'h00000000 /* 0xb48c */;
                11556: data_o = 32'h00000000 /* 0xb490 */;
                11557: data_o = 32'h00000000 /* 0xb494 */;
                11558: data_o = 32'h00000000 /* 0xb498 */;
                11559: data_o = 32'h00000000 /* 0xb49c */;
                11560: data_o = 32'h00000000 /* 0xb4a0 */;
                11561: data_o = 32'h00000000 /* 0xb4a4 */;
                11562: data_o = 32'h00000000 /* 0xb4a8 */;
                11563: data_o = 32'h00000000 /* 0xb4ac */;
                11564: data_o = 32'h00000000 /* 0xb4b0 */;
                11565: data_o = 32'h00000000 /* 0xb4b4 */;
                11566: data_o = 32'h00000000 /* 0xb4b8 */;
                11567: data_o = 32'h00000000 /* 0xb4bc */;
                11568: data_o = 32'h00000000 /* 0xb4c0 */;
                11569: data_o = 32'h00000000 /* 0xb4c4 */;
                11570: data_o = 32'h00000000 /* 0xb4c8 */;
                11571: data_o = 32'h00000000 /* 0xb4cc */;
                11572: data_o = 32'h00000000 /* 0xb4d0 */;
                11573: data_o = 32'h00000000 /* 0xb4d4 */;
                11574: data_o = 32'h00000000 /* 0xb4d8 */;
                11575: data_o = 32'h00000000 /* 0xb4dc */;
                11576: data_o = 32'h00000000 /* 0xb4e0 */;
                11577: data_o = 32'h00000000 /* 0xb4e4 */;
                11578: data_o = 32'h00000000 /* 0xb4e8 */;
                11579: data_o = 32'h00000000 /* 0xb4ec */;
                11580: data_o = 32'h00000000 /* 0xb4f0 */;
                11581: data_o = 32'h00000000 /* 0xb4f4 */;
                11582: data_o = 32'h00000000 /* 0xb4f8 */;
                11583: data_o = 32'h00000000 /* 0xb4fc */;
                11584: data_o = 32'h00000000 /* 0xb500 */;
                11585: data_o = 32'h00000000 /* 0xb504 */;
                11586: data_o = 32'h00000000 /* 0xb508 */;
                11587: data_o = 32'h00000000 /* 0xb50c */;
                11588: data_o = 32'h00000000 /* 0xb510 */;
                11589: data_o = 32'h00000000 /* 0xb514 */;
                11590: data_o = 32'h00000000 /* 0xb518 */;
                11591: data_o = 32'h00000000 /* 0xb51c */;
                11592: data_o = 32'h00000000 /* 0xb520 */;
                11593: data_o = 32'h00000000 /* 0xb524 */;
                11594: data_o = 32'h00000000 /* 0xb528 */;
                11595: data_o = 32'h00000000 /* 0xb52c */;
                11596: data_o = 32'h00000000 /* 0xb530 */;
                11597: data_o = 32'h00000000 /* 0xb534 */;
                11598: data_o = 32'h00000000 /* 0xb538 */;
                11599: data_o = 32'h00000000 /* 0xb53c */;
                11600: data_o = 32'h00000000 /* 0xb540 */;
                11601: data_o = 32'h00000000 /* 0xb544 */;
                11602: data_o = 32'h00000000 /* 0xb548 */;
                11603: data_o = 32'h00000000 /* 0xb54c */;
                11604: data_o = 32'h00000000 /* 0xb550 */;
                11605: data_o = 32'h00000000 /* 0xb554 */;
                11606: data_o = 32'h00000000 /* 0xb558 */;
                11607: data_o = 32'h00000000 /* 0xb55c */;
                11608: data_o = 32'h00000000 /* 0xb560 */;
                11609: data_o = 32'h00000000 /* 0xb564 */;
                11610: data_o = 32'h00000000 /* 0xb568 */;
                11611: data_o = 32'h00000000 /* 0xb56c */;
                11612: data_o = 32'h00000000 /* 0xb570 */;
                11613: data_o = 32'h00000000 /* 0xb574 */;
                11614: data_o = 32'h00000000 /* 0xb578 */;
                11615: data_o = 32'h00000000 /* 0xb57c */;
                11616: data_o = 32'h00000000 /* 0xb580 */;
                11617: data_o = 32'h00000000 /* 0xb584 */;
                11618: data_o = 32'h00000000 /* 0xb588 */;
                11619: data_o = 32'h00000000 /* 0xb58c */;
                11620: data_o = 32'h00000000 /* 0xb590 */;
                11621: data_o = 32'h00000000 /* 0xb594 */;
                11622: data_o = 32'h00000000 /* 0xb598 */;
                11623: data_o = 32'h00000000 /* 0xb59c */;
                11624: data_o = 32'h00000000 /* 0xb5a0 */;
                11625: data_o = 32'h00000000 /* 0xb5a4 */;
                11626: data_o = 32'h00000000 /* 0xb5a8 */;
                11627: data_o = 32'h00000000 /* 0xb5ac */;
                11628: data_o = 32'h00000000 /* 0xb5b0 */;
                11629: data_o = 32'h00000000 /* 0xb5b4 */;
                11630: data_o = 32'h00000000 /* 0xb5b8 */;
                11631: data_o = 32'h00000000 /* 0xb5bc */;
                11632: data_o = 32'h00000000 /* 0xb5c0 */;
                11633: data_o = 32'h00000000 /* 0xb5c4 */;
                11634: data_o = 32'h00000000 /* 0xb5c8 */;
                11635: data_o = 32'h00000000 /* 0xb5cc */;
                11636: data_o = 32'h00000000 /* 0xb5d0 */;
                11637: data_o = 32'h00000000 /* 0xb5d4 */;
                11638: data_o = 32'h00000000 /* 0xb5d8 */;
                11639: data_o = 32'h00000000 /* 0xb5dc */;
                11640: data_o = 32'h00000000 /* 0xb5e0 */;
                11641: data_o = 32'h00000000 /* 0xb5e4 */;
                11642: data_o = 32'h00000000 /* 0xb5e8 */;
                11643: data_o = 32'h00000000 /* 0xb5ec */;
                11644: data_o = 32'h00000000 /* 0xb5f0 */;
                11645: data_o = 32'h00000000 /* 0xb5f4 */;
                11646: data_o = 32'h00000000 /* 0xb5f8 */;
                11647: data_o = 32'h00000000 /* 0xb5fc */;
                11648: data_o = 32'h00000000 /* 0xb600 */;
                11649: data_o = 32'h00000000 /* 0xb604 */;
                11650: data_o = 32'h00000000 /* 0xb608 */;
                11651: data_o = 32'h00000000 /* 0xb60c */;
                11652: data_o = 32'h00000000 /* 0xb610 */;
                11653: data_o = 32'h00000000 /* 0xb614 */;
                11654: data_o = 32'h00000000 /* 0xb618 */;
                11655: data_o = 32'h00000000 /* 0xb61c */;
                11656: data_o = 32'h00000000 /* 0xb620 */;
                11657: data_o = 32'h00000000 /* 0xb624 */;
                11658: data_o = 32'h00000000 /* 0xb628 */;
                11659: data_o = 32'h00000000 /* 0xb62c */;
                11660: data_o = 32'h00000000 /* 0xb630 */;
                11661: data_o = 32'h00000000 /* 0xb634 */;
                11662: data_o = 32'h00000000 /* 0xb638 */;
                11663: data_o = 32'h00000000 /* 0xb63c */;
                11664: data_o = 32'h00000000 /* 0xb640 */;
                11665: data_o = 32'h00000000 /* 0xb644 */;
                11666: data_o = 32'h00000000 /* 0xb648 */;
                11667: data_o = 32'h00000000 /* 0xb64c */;
                11668: data_o = 32'h00000000 /* 0xb650 */;
                11669: data_o = 32'h00000000 /* 0xb654 */;
                11670: data_o = 32'h00000000 /* 0xb658 */;
                11671: data_o = 32'h00000000 /* 0xb65c */;
                11672: data_o = 32'h00000000 /* 0xb660 */;
                11673: data_o = 32'h00000000 /* 0xb664 */;
                11674: data_o = 32'h00000000 /* 0xb668 */;
                11675: data_o = 32'h00000000 /* 0xb66c */;
                11676: data_o = 32'h00000000 /* 0xb670 */;
                11677: data_o = 32'h00000000 /* 0xb674 */;
                11678: data_o = 32'h00000000 /* 0xb678 */;
                11679: data_o = 32'h00000000 /* 0xb67c */;
                11680: data_o = 32'h00000000 /* 0xb680 */;
                11681: data_o = 32'h00000000 /* 0xb684 */;
                11682: data_o = 32'h00000000 /* 0xb688 */;
                11683: data_o = 32'h00000000 /* 0xb68c */;
                11684: data_o = 32'h00000000 /* 0xb690 */;
                11685: data_o = 32'h00000000 /* 0xb694 */;
                11686: data_o = 32'h00000000 /* 0xb698 */;
                11687: data_o = 32'h00000000 /* 0xb69c */;
                11688: data_o = 32'h00000000 /* 0xb6a0 */;
                11689: data_o = 32'h00000000 /* 0xb6a4 */;
                11690: data_o = 32'h00000000 /* 0xb6a8 */;
                11691: data_o = 32'h00000000 /* 0xb6ac */;
                11692: data_o = 32'h00000000 /* 0xb6b0 */;
                11693: data_o = 32'h00000000 /* 0xb6b4 */;
                11694: data_o = 32'h00000000 /* 0xb6b8 */;
                11695: data_o = 32'h00000000 /* 0xb6bc */;
                11696: data_o = 32'h00000000 /* 0xb6c0 */;
                11697: data_o = 32'h00000000 /* 0xb6c4 */;
                11698: data_o = 32'h00000000 /* 0xb6c8 */;
                11699: data_o = 32'h00000000 /* 0xb6cc */;
                11700: data_o = 32'h00000000 /* 0xb6d0 */;
                11701: data_o = 32'h00000000 /* 0xb6d4 */;
                11702: data_o = 32'h00000000 /* 0xb6d8 */;
                11703: data_o = 32'h00000000 /* 0xb6dc */;
                11704: data_o = 32'h00000000 /* 0xb6e0 */;
                11705: data_o = 32'h00000000 /* 0xb6e4 */;
                11706: data_o = 32'h00000000 /* 0xb6e8 */;
                11707: data_o = 32'h00000000 /* 0xb6ec */;
                11708: data_o = 32'h00000000 /* 0xb6f0 */;
                11709: data_o = 32'h00000000 /* 0xb6f4 */;
                11710: data_o = 32'h00000000 /* 0xb6f8 */;
                11711: data_o = 32'h00000000 /* 0xb6fc */;
                11712: data_o = 32'h00000000 /* 0xb700 */;
                11713: data_o = 32'h00000000 /* 0xb704 */;
                11714: data_o = 32'h00000000 /* 0xb708 */;
                11715: data_o = 32'h00000000 /* 0xb70c */;
                11716: data_o = 32'h00000000 /* 0xb710 */;
                11717: data_o = 32'h00000000 /* 0xb714 */;
                11718: data_o = 32'h00000000 /* 0xb718 */;
                11719: data_o = 32'h00000000 /* 0xb71c */;
                11720: data_o = 32'h00000000 /* 0xb720 */;
                11721: data_o = 32'h00000000 /* 0xb724 */;
                11722: data_o = 32'h00000000 /* 0xb728 */;
                11723: data_o = 32'h00000000 /* 0xb72c */;
                11724: data_o = 32'h00000000 /* 0xb730 */;
                11725: data_o = 32'h00000000 /* 0xb734 */;
                11726: data_o = 32'h00000000 /* 0xb738 */;
                11727: data_o = 32'h00000000 /* 0xb73c */;
                11728: data_o = 32'h00000000 /* 0xb740 */;
                11729: data_o = 32'h00000000 /* 0xb744 */;
                11730: data_o = 32'h00000000 /* 0xb748 */;
                11731: data_o = 32'h00000000 /* 0xb74c */;
                11732: data_o = 32'h00000000 /* 0xb750 */;
                11733: data_o = 32'h00000000 /* 0xb754 */;
                11734: data_o = 32'h00000000 /* 0xb758 */;
                11735: data_o = 32'h00000000 /* 0xb75c */;
                11736: data_o = 32'h00000000 /* 0xb760 */;
                11737: data_o = 32'h00000000 /* 0xb764 */;
                11738: data_o = 32'h00000000 /* 0xb768 */;
                11739: data_o = 32'h00000000 /* 0xb76c */;
                11740: data_o = 32'h00000000 /* 0xb770 */;
                11741: data_o = 32'h00000000 /* 0xb774 */;
                11742: data_o = 32'h00000000 /* 0xb778 */;
                11743: data_o = 32'h00000000 /* 0xb77c */;
                11744: data_o = 32'h00000000 /* 0xb780 */;
                11745: data_o = 32'h00000000 /* 0xb784 */;
                11746: data_o = 32'h00000000 /* 0xb788 */;
                11747: data_o = 32'h00000000 /* 0xb78c */;
                11748: data_o = 32'h00000000 /* 0xb790 */;
                11749: data_o = 32'h00000000 /* 0xb794 */;
                11750: data_o = 32'h00000000 /* 0xb798 */;
                11751: data_o = 32'h00000000 /* 0xb79c */;
                11752: data_o = 32'h00000000 /* 0xb7a0 */;
                11753: data_o = 32'h00000000 /* 0xb7a4 */;
                11754: data_o = 32'h00000000 /* 0xb7a8 */;
                11755: data_o = 32'h00000000 /* 0xb7ac */;
                11756: data_o = 32'h00000000 /* 0xb7b0 */;
                11757: data_o = 32'h00000000 /* 0xb7b4 */;
                11758: data_o = 32'h00000000 /* 0xb7b8 */;
                11759: data_o = 32'h00000000 /* 0xb7bc */;
                11760: data_o = 32'h00000000 /* 0xb7c0 */;
                11761: data_o = 32'h00000000 /* 0xb7c4 */;
                11762: data_o = 32'h00000000 /* 0xb7c8 */;
                11763: data_o = 32'h00000000 /* 0xb7cc */;
                11764: data_o = 32'h00000000 /* 0xb7d0 */;
                11765: data_o = 32'h00000000 /* 0xb7d4 */;
                11766: data_o = 32'h00000000 /* 0xb7d8 */;
                11767: data_o = 32'h00000000 /* 0xb7dc */;
                11768: data_o = 32'h00000000 /* 0xb7e0 */;
                11769: data_o = 32'h00000000 /* 0xb7e4 */;
                11770: data_o = 32'h00000000 /* 0xb7e8 */;
                11771: data_o = 32'h00000000 /* 0xb7ec */;
                11772: data_o = 32'h00000000 /* 0xb7f0 */;
                11773: data_o = 32'h00000000 /* 0xb7f4 */;
                11774: data_o = 32'h00000000 /* 0xb7f8 */;
                11775: data_o = 32'h00000000 /* 0xb7fc */;
                11776: data_o = 32'h00000000 /* 0xb800 */;
                11777: data_o = 32'h00000000 /* 0xb804 */;
                11778: data_o = 32'h00000000 /* 0xb808 */;
                11779: data_o = 32'h00000000 /* 0xb80c */;
                11780: data_o = 32'h00000000 /* 0xb810 */;
                11781: data_o = 32'h00000000 /* 0xb814 */;
                11782: data_o = 32'h00000000 /* 0xb818 */;
                11783: data_o = 32'h00000000 /* 0xb81c */;
                11784: data_o = 32'h00000000 /* 0xb820 */;
                11785: data_o = 32'h00000000 /* 0xb824 */;
                11786: data_o = 32'h00000000 /* 0xb828 */;
                11787: data_o = 32'h00000000 /* 0xb82c */;
                11788: data_o = 32'h00000000 /* 0xb830 */;
                11789: data_o = 32'h00000000 /* 0xb834 */;
                11790: data_o = 32'h00000000 /* 0xb838 */;
                11791: data_o = 32'h00000000 /* 0xb83c */;
                11792: data_o = 32'h00000000 /* 0xb840 */;
                11793: data_o = 32'h00000000 /* 0xb844 */;
                11794: data_o = 32'h00000000 /* 0xb848 */;
                11795: data_o = 32'h00000000 /* 0xb84c */;
                11796: data_o = 32'h00000000 /* 0xb850 */;
                11797: data_o = 32'h00000000 /* 0xb854 */;
                11798: data_o = 32'h00000000 /* 0xb858 */;
                11799: data_o = 32'h00000000 /* 0xb85c */;
                11800: data_o = 32'h00000000 /* 0xb860 */;
                11801: data_o = 32'h00000000 /* 0xb864 */;
                11802: data_o = 32'h00000000 /* 0xb868 */;
                11803: data_o = 32'h00000000 /* 0xb86c */;
                11804: data_o = 32'h00000000 /* 0xb870 */;
                11805: data_o = 32'h00000000 /* 0xb874 */;
                11806: data_o = 32'h00000000 /* 0xb878 */;
                11807: data_o = 32'h00000000 /* 0xb87c */;
                11808: data_o = 32'h00000000 /* 0xb880 */;
                11809: data_o = 32'h00000000 /* 0xb884 */;
                11810: data_o = 32'h00000000 /* 0xb888 */;
                11811: data_o = 32'h00000000 /* 0xb88c */;
                11812: data_o = 32'h00000000 /* 0xb890 */;
                11813: data_o = 32'h00000000 /* 0xb894 */;
                11814: data_o = 32'h00000000 /* 0xb898 */;
                11815: data_o = 32'h00000000 /* 0xb89c */;
                11816: data_o = 32'h00000000 /* 0xb8a0 */;
                11817: data_o = 32'h00000000 /* 0xb8a4 */;
                11818: data_o = 32'h00000000 /* 0xb8a8 */;
                11819: data_o = 32'h00000000 /* 0xb8ac */;
                11820: data_o = 32'h00000000 /* 0xb8b0 */;
                11821: data_o = 32'h00000000 /* 0xb8b4 */;
                11822: data_o = 32'h00000000 /* 0xb8b8 */;
                11823: data_o = 32'h00000000 /* 0xb8bc */;
                11824: data_o = 32'h00000000 /* 0xb8c0 */;
                11825: data_o = 32'h00000000 /* 0xb8c4 */;
                11826: data_o = 32'h00000000 /* 0xb8c8 */;
                11827: data_o = 32'h00000000 /* 0xb8cc */;
                11828: data_o = 32'h00000000 /* 0xb8d0 */;
                11829: data_o = 32'h00000000 /* 0xb8d4 */;
                11830: data_o = 32'h00000000 /* 0xb8d8 */;
                11831: data_o = 32'h00000000 /* 0xb8dc */;
                11832: data_o = 32'h00000000 /* 0xb8e0 */;
                11833: data_o = 32'h00000000 /* 0xb8e4 */;
                11834: data_o = 32'h00000000 /* 0xb8e8 */;
                11835: data_o = 32'h00000000 /* 0xb8ec */;
                11836: data_o = 32'h00000000 /* 0xb8f0 */;
                11837: data_o = 32'h00000000 /* 0xb8f4 */;
                11838: data_o = 32'h00000000 /* 0xb8f8 */;
                11839: data_o = 32'h00000000 /* 0xb8fc */;
                11840: data_o = 32'h00000000 /* 0xb900 */;
                11841: data_o = 32'h00000000 /* 0xb904 */;
                11842: data_o = 32'h00000000 /* 0xb908 */;
                11843: data_o = 32'h00000000 /* 0xb90c */;
                11844: data_o = 32'h00000000 /* 0xb910 */;
                11845: data_o = 32'h00000000 /* 0xb914 */;
                11846: data_o = 32'h00000000 /* 0xb918 */;
                11847: data_o = 32'h00000000 /* 0xb91c */;
                11848: data_o = 32'h00000000 /* 0xb920 */;
                11849: data_o = 32'h00000000 /* 0xb924 */;
                11850: data_o = 32'h00000000 /* 0xb928 */;
                11851: data_o = 32'h00000000 /* 0xb92c */;
                11852: data_o = 32'h00000000 /* 0xb930 */;
                11853: data_o = 32'h00000000 /* 0xb934 */;
                11854: data_o = 32'h00000000 /* 0xb938 */;
                11855: data_o = 32'h00000000 /* 0xb93c */;
                11856: data_o = 32'h00000000 /* 0xb940 */;
                11857: data_o = 32'h00000000 /* 0xb944 */;
                11858: data_o = 32'h00000000 /* 0xb948 */;
                11859: data_o = 32'h00000000 /* 0xb94c */;
                11860: data_o = 32'h00000000 /* 0xb950 */;
                11861: data_o = 32'h00000000 /* 0xb954 */;
                11862: data_o = 32'h00000000 /* 0xb958 */;
                11863: data_o = 32'h00000000 /* 0xb95c */;
                11864: data_o = 32'h00000000 /* 0xb960 */;
                11865: data_o = 32'h00000000 /* 0xb964 */;
                11866: data_o = 32'h00000000 /* 0xb968 */;
                11867: data_o = 32'h00000000 /* 0xb96c */;
                11868: data_o = 32'h00000000 /* 0xb970 */;
                11869: data_o = 32'h00000000 /* 0xb974 */;
                11870: data_o = 32'h00000000 /* 0xb978 */;
                11871: data_o = 32'h00000000 /* 0xb97c */;
                11872: data_o = 32'h00000000 /* 0xb980 */;
                11873: data_o = 32'h00000000 /* 0xb984 */;
                11874: data_o = 32'h00000000 /* 0xb988 */;
                11875: data_o = 32'h00000000 /* 0xb98c */;
                11876: data_o = 32'h00000000 /* 0xb990 */;
                11877: data_o = 32'h00000000 /* 0xb994 */;
                11878: data_o = 32'h00000000 /* 0xb998 */;
                11879: data_o = 32'h00000000 /* 0xb99c */;
                11880: data_o = 32'h00000000 /* 0xb9a0 */;
                11881: data_o = 32'h00000000 /* 0xb9a4 */;
                11882: data_o = 32'h00000000 /* 0xb9a8 */;
                11883: data_o = 32'h00000000 /* 0xb9ac */;
                11884: data_o = 32'h00000000 /* 0xb9b0 */;
                11885: data_o = 32'h00000000 /* 0xb9b4 */;
                11886: data_o = 32'h00000000 /* 0xb9b8 */;
                11887: data_o = 32'h00000000 /* 0xb9bc */;
                11888: data_o = 32'h00000000 /* 0xb9c0 */;
                11889: data_o = 32'h00000000 /* 0xb9c4 */;
                11890: data_o = 32'h00000000 /* 0xb9c8 */;
                11891: data_o = 32'h00000000 /* 0xb9cc */;
                11892: data_o = 32'h00000000 /* 0xb9d0 */;
                11893: data_o = 32'h00000000 /* 0xb9d4 */;
                11894: data_o = 32'h00000000 /* 0xb9d8 */;
                11895: data_o = 32'h00000000 /* 0xb9dc */;
                11896: data_o = 32'h00000000 /* 0xb9e0 */;
                11897: data_o = 32'h00000000 /* 0xb9e4 */;
                11898: data_o = 32'h00000000 /* 0xb9e8 */;
                11899: data_o = 32'h00000000 /* 0xb9ec */;
                11900: data_o = 32'h00000000 /* 0xb9f0 */;
                11901: data_o = 32'h00000000 /* 0xb9f4 */;
                11902: data_o = 32'h00000000 /* 0xb9f8 */;
                11903: data_o = 32'h00000000 /* 0xb9fc */;
                11904: data_o = 32'h00000000 /* 0xba00 */;
                11905: data_o = 32'h00000000 /* 0xba04 */;
                11906: data_o = 32'h00000000 /* 0xba08 */;
                11907: data_o = 32'h00000000 /* 0xba0c */;
                11908: data_o = 32'h00000000 /* 0xba10 */;
                11909: data_o = 32'h00000000 /* 0xba14 */;
                11910: data_o = 32'h00000000 /* 0xba18 */;
                11911: data_o = 32'h00000000 /* 0xba1c */;
                11912: data_o = 32'h00000000 /* 0xba20 */;
                11913: data_o = 32'h00000000 /* 0xba24 */;
                11914: data_o = 32'h00000000 /* 0xba28 */;
                11915: data_o = 32'h00000000 /* 0xba2c */;
                11916: data_o = 32'h00000000 /* 0xba30 */;
                11917: data_o = 32'h00000000 /* 0xba34 */;
                11918: data_o = 32'h00000000 /* 0xba38 */;
                11919: data_o = 32'h00000000 /* 0xba3c */;
                11920: data_o = 32'h00000000 /* 0xba40 */;
                11921: data_o = 32'h00000000 /* 0xba44 */;
                11922: data_o = 32'h00000000 /* 0xba48 */;
                11923: data_o = 32'h00000000 /* 0xba4c */;
                11924: data_o = 32'h00000000 /* 0xba50 */;
                11925: data_o = 32'h00000000 /* 0xba54 */;
                11926: data_o = 32'h00000000 /* 0xba58 */;
                11927: data_o = 32'h00000000 /* 0xba5c */;
                11928: data_o = 32'h00000000 /* 0xba60 */;
                11929: data_o = 32'h00000000 /* 0xba64 */;
                11930: data_o = 32'h00000000 /* 0xba68 */;
                11931: data_o = 32'h00000000 /* 0xba6c */;
                11932: data_o = 32'h00000000 /* 0xba70 */;
                11933: data_o = 32'h00000000 /* 0xba74 */;
                11934: data_o = 32'h00000000 /* 0xba78 */;
                11935: data_o = 32'h00000000 /* 0xba7c */;
                11936: data_o = 32'h00000000 /* 0xba80 */;
                11937: data_o = 32'h00000000 /* 0xba84 */;
                11938: data_o = 32'h00000000 /* 0xba88 */;
                11939: data_o = 32'h00000000 /* 0xba8c */;
                11940: data_o = 32'h00000000 /* 0xba90 */;
                11941: data_o = 32'h00000000 /* 0xba94 */;
                11942: data_o = 32'h00000000 /* 0xba98 */;
                11943: data_o = 32'h00000000 /* 0xba9c */;
                11944: data_o = 32'h00000000 /* 0xbaa0 */;
                11945: data_o = 32'h00000000 /* 0xbaa4 */;
                11946: data_o = 32'h00000000 /* 0xbaa8 */;
                11947: data_o = 32'h00000000 /* 0xbaac */;
                11948: data_o = 32'h00000000 /* 0xbab0 */;
                11949: data_o = 32'h00000000 /* 0xbab4 */;
                11950: data_o = 32'h00000000 /* 0xbab8 */;
                11951: data_o = 32'h00000000 /* 0xbabc */;
                11952: data_o = 32'h00000000 /* 0xbac0 */;
                11953: data_o = 32'h00000000 /* 0xbac4 */;
                11954: data_o = 32'h00000000 /* 0xbac8 */;
                11955: data_o = 32'h00000000 /* 0xbacc */;
                11956: data_o = 32'h00000000 /* 0xbad0 */;
                11957: data_o = 32'h00000000 /* 0xbad4 */;
                11958: data_o = 32'h00000000 /* 0xbad8 */;
                11959: data_o = 32'h00000000 /* 0xbadc */;
                11960: data_o = 32'h00000000 /* 0xbae0 */;
                11961: data_o = 32'h00000000 /* 0xbae4 */;
                11962: data_o = 32'h00000000 /* 0xbae8 */;
                11963: data_o = 32'h00000000 /* 0xbaec */;
                11964: data_o = 32'h00000000 /* 0xbaf0 */;
                11965: data_o = 32'h00000000 /* 0xbaf4 */;
                11966: data_o = 32'h00000000 /* 0xbaf8 */;
                11967: data_o = 32'h00000000 /* 0xbafc */;
                11968: data_o = 32'h00000000 /* 0xbb00 */;
                11969: data_o = 32'h00000000 /* 0xbb04 */;
                11970: data_o = 32'h00000000 /* 0xbb08 */;
                11971: data_o = 32'h00000000 /* 0xbb0c */;
                11972: data_o = 32'h00000000 /* 0xbb10 */;
                11973: data_o = 32'h00000000 /* 0xbb14 */;
                11974: data_o = 32'h00000000 /* 0xbb18 */;
                11975: data_o = 32'h00000000 /* 0xbb1c */;
                11976: data_o = 32'h00000000 /* 0xbb20 */;
                11977: data_o = 32'h00000000 /* 0xbb24 */;
                11978: data_o = 32'h00000000 /* 0xbb28 */;
                11979: data_o = 32'h00000000 /* 0xbb2c */;
                11980: data_o = 32'h00000000 /* 0xbb30 */;
                11981: data_o = 32'h00000000 /* 0xbb34 */;
                11982: data_o = 32'h00000000 /* 0xbb38 */;
                11983: data_o = 32'h00000000 /* 0xbb3c */;
                11984: data_o = 32'h00000000 /* 0xbb40 */;
                11985: data_o = 32'h00000000 /* 0xbb44 */;
                11986: data_o = 32'h00000000 /* 0xbb48 */;
                11987: data_o = 32'h00000000 /* 0xbb4c */;
                11988: data_o = 32'h00000000 /* 0xbb50 */;
                11989: data_o = 32'h00000000 /* 0xbb54 */;
                11990: data_o = 32'h00000000 /* 0xbb58 */;
                11991: data_o = 32'h00000000 /* 0xbb5c */;
                11992: data_o = 32'h00000000 /* 0xbb60 */;
                11993: data_o = 32'h00000000 /* 0xbb64 */;
                11994: data_o = 32'h00000000 /* 0xbb68 */;
                11995: data_o = 32'h00000000 /* 0xbb6c */;
                11996: data_o = 32'h00000000 /* 0xbb70 */;
                11997: data_o = 32'h00000000 /* 0xbb74 */;
                11998: data_o = 32'h00000000 /* 0xbb78 */;
                11999: data_o = 32'h00000000 /* 0xbb7c */;
                12000: data_o = 32'h00000000 /* 0xbb80 */;
                12001: data_o = 32'h00000000 /* 0xbb84 */;
                12002: data_o = 32'h00000000 /* 0xbb88 */;
                12003: data_o = 32'h00000000 /* 0xbb8c */;
                12004: data_o = 32'h00000000 /* 0xbb90 */;
                12005: data_o = 32'h00000000 /* 0xbb94 */;
                12006: data_o = 32'h00000000 /* 0xbb98 */;
                12007: data_o = 32'h00000000 /* 0xbb9c */;
                12008: data_o = 32'h00000000 /* 0xbba0 */;
                12009: data_o = 32'h00000000 /* 0xbba4 */;
                12010: data_o = 32'h00000000 /* 0xbba8 */;
                12011: data_o = 32'h00000000 /* 0xbbac */;
                12012: data_o = 32'h00000000 /* 0xbbb0 */;
                12013: data_o = 32'h00000000 /* 0xbbb4 */;
                12014: data_o = 32'h00000000 /* 0xbbb8 */;
                12015: data_o = 32'h00000000 /* 0xbbbc */;
                12016: data_o = 32'h00000000 /* 0xbbc0 */;
                12017: data_o = 32'h00000000 /* 0xbbc4 */;
                12018: data_o = 32'h00000000 /* 0xbbc8 */;
                12019: data_o = 32'h00000000 /* 0xbbcc */;
                12020: data_o = 32'h00000000 /* 0xbbd0 */;
                12021: data_o = 32'h00000000 /* 0xbbd4 */;
                12022: data_o = 32'h00000000 /* 0xbbd8 */;
                12023: data_o = 32'h00000000 /* 0xbbdc */;
                12024: data_o = 32'h00000000 /* 0xbbe0 */;
                12025: data_o = 32'h00000000 /* 0xbbe4 */;
                12026: data_o = 32'h00000000 /* 0xbbe8 */;
                12027: data_o = 32'h00000000 /* 0xbbec */;
                12028: data_o = 32'h00000000 /* 0xbbf0 */;
                12029: data_o = 32'h00000000 /* 0xbbf4 */;
                12030: data_o = 32'h00000000 /* 0xbbf8 */;
                12031: data_o = 32'h00000000 /* 0xbbfc */;
                12032: data_o = 32'h00000000 /* 0xbc00 */;
                12033: data_o = 32'h00000000 /* 0xbc04 */;
                12034: data_o = 32'h00000000 /* 0xbc08 */;
                12035: data_o = 32'h00000000 /* 0xbc0c */;
                12036: data_o = 32'h00000000 /* 0xbc10 */;
                12037: data_o = 32'h00000000 /* 0xbc14 */;
                12038: data_o = 32'h00000000 /* 0xbc18 */;
                12039: data_o = 32'h00000000 /* 0xbc1c */;
                12040: data_o = 32'h00000000 /* 0xbc20 */;
                12041: data_o = 32'h00000000 /* 0xbc24 */;
                12042: data_o = 32'h00000000 /* 0xbc28 */;
                12043: data_o = 32'h00000000 /* 0xbc2c */;
                12044: data_o = 32'h00000000 /* 0xbc30 */;
                12045: data_o = 32'h00000000 /* 0xbc34 */;
                12046: data_o = 32'h00000000 /* 0xbc38 */;
                12047: data_o = 32'h00000000 /* 0xbc3c */;
                12048: data_o = 32'h00000000 /* 0xbc40 */;
                12049: data_o = 32'h00000000 /* 0xbc44 */;
                12050: data_o = 32'h00000000 /* 0xbc48 */;
                12051: data_o = 32'h00000000 /* 0xbc4c */;
                12052: data_o = 32'h00000000 /* 0xbc50 */;
                12053: data_o = 32'h00000000 /* 0xbc54 */;
                12054: data_o = 32'h00000000 /* 0xbc58 */;
                12055: data_o = 32'h00000000 /* 0xbc5c */;
                12056: data_o = 32'h00000000 /* 0xbc60 */;
                12057: data_o = 32'h00000000 /* 0xbc64 */;
                12058: data_o = 32'h00000000 /* 0xbc68 */;
                12059: data_o = 32'h00000000 /* 0xbc6c */;
                12060: data_o = 32'h00000000 /* 0xbc70 */;
                12061: data_o = 32'h00000000 /* 0xbc74 */;
                12062: data_o = 32'h00000000 /* 0xbc78 */;
                12063: data_o = 32'h00000000 /* 0xbc7c */;
                12064: data_o = 32'h00000000 /* 0xbc80 */;
                12065: data_o = 32'h00000000 /* 0xbc84 */;
                12066: data_o = 32'h00000000 /* 0xbc88 */;
                12067: data_o = 32'h00000000 /* 0xbc8c */;
                12068: data_o = 32'h00000000 /* 0xbc90 */;
                12069: data_o = 32'h00000000 /* 0xbc94 */;
                12070: data_o = 32'h00000000 /* 0xbc98 */;
                12071: data_o = 32'h00000000 /* 0xbc9c */;
                12072: data_o = 32'h00000000 /* 0xbca0 */;
                12073: data_o = 32'h00000000 /* 0xbca4 */;
                12074: data_o = 32'h00000000 /* 0xbca8 */;
                12075: data_o = 32'h00000000 /* 0xbcac */;
                12076: data_o = 32'h00000000 /* 0xbcb0 */;
                12077: data_o = 32'h00000000 /* 0xbcb4 */;
                12078: data_o = 32'h00000000 /* 0xbcb8 */;
                12079: data_o = 32'h00000000 /* 0xbcbc */;
                12080: data_o = 32'h00000000 /* 0xbcc0 */;
                12081: data_o = 32'h00000000 /* 0xbcc4 */;
                12082: data_o = 32'h00000000 /* 0xbcc8 */;
                12083: data_o = 32'h00000000 /* 0xbccc */;
                12084: data_o = 32'h00000000 /* 0xbcd0 */;
                12085: data_o = 32'h00000000 /* 0xbcd4 */;
                12086: data_o = 32'h00000000 /* 0xbcd8 */;
                12087: data_o = 32'h00000000 /* 0xbcdc */;
                12088: data_o = 32'h00000000 /* 0xbce0 */;
                12089: data_o = 32'h00000000 /* 0xbce4 */;
                12090: data_o = 32'h00000000 /* 0xbce8 */;
                12091: data_o = 32'h00000000 /* 0xbcec */;
                12092: data_o = 32'h00000000 /* 0xbcf0 */;
                12093: data_o = 32'h00000000 /* 0xbcf4 */;
                12094: data_o = 32'h00000000 /* 0xbcf8 */;
                12095: data_o = 32'h00000000 /* 0xbcfc */;
                12096: data_o = 32'h00000000 /* 0xbd00 */;
                12097: data_o = 32'h00000000 /* 0xbd04 */;
                12098: data_o = 32'h00000000 /* 0xbd08 */;
                12099: data_o = 32'h00000000 /* 0xbd0c */;
                12100: data_o = 32'h00000000 /* 0xbd10 */;
                12101: data_o = 32'h00000000 /* 0xbd14 */;
                12102: data_o = 32'h00000000 /* 0xbd18 */;
                12103: data_o = 32'h00000000 /* 0xbd1c */;
                12104: data_o = 32'h00000000 /* 0xbd20 */;
                12105: data_o = 32'h00000000 /* 0xbd24 */;
                12106: data_o = 32'h00000000 /* 0xbd28 */;
                12107: data_o = 32'h00000000 /* 0xbd2c */;
                12108: data_o = 32'h00000000 /* 0xbd30 */;
                12109: data_o = 32'h00000000 /* 0xbd34 */;
                12110: data_o = 32'h00000000 /* 0xbd38 */;
                12111: data_o = 32'h00000000 /* 0xbd3c */;
                12112: data_o = 32'h00000000 /* 0xbd40 */;
                12113: data_o = 32'h00000000 /* 0xbd44 */;
                12114: data_o = 32'h00000000 /* 0xbd48 */;
                12115: data_o = 32'h00000000 /* 0xbd4c */;
                12116: data_o = 32'h00000000 /* 0xbd50 */;
                12117: data_o = 32'h00000000 /* 0xbd54 */;
                12118: data_o = 32'h00000000 /* 0xbd58 */;
                12119: data_o = 32'h00000000 /* 0xbd5c */;
                12120: data_o = 32'h00000000 /* 0xbd60 */;
                12121: data_o = 32'h00000000 /* 0xbd64 */;
                12122: data_o = 32'h00000000 /* 0xbd68 */;
                12123: data_o = 32'h00000000 /* 0xbd6c */;
                12124: data_o = 32'h00000000 /* 0xbd70 */;
                12125: data_o = 32'h00000000 /* 0xbd74 */;
                12126: data_o = 32'h00000000 /* 0xbd78 */;
                12127: data_o = 32'h00000000 /* 0xbd7c */;
                12128: data_o = 32'h00000000 /* 0xbd80 */;
                12129: data_o = 32'h00000000 /* 0xbd84 */;
                12130: data_o = 32'h00000000 /* 0xbd88 */;
                12131: data_o = 32'h00000000 /* 0xbd8c */;
                12132: data_o = 32'h00000000 /* 0xbd90 */;
                12133: data_o = 32'h00000000 /* 0xbd94 */;
                12134: data_o = 32'h00000000 /* 0xbd98 */;
                12135: data_o = 32'h00000000 /* 0xbd9c */;
                12136: data_o = 32'h00000000 /* 0xbda0 */;
                12137: data_o = 32'h00000000 /* 0xbda4 */;
                12138: data_o = 32'h00000000 /* 0xbda8 */;
                12139: data_o = 32'h00000000 /* 0xbdac */;
                12140: data_o = 32'h00000000 /* 0xbdb0 */;
                12141: data_o = 32'h00000000 /* 0xbdb4 */;
                12142: data_o = 32'h00000000 /* 0xbdb8 */;
                12143: data_o = 32'h00000000 /* 0xbdbc */;
                12144: data_o = 32'h00000000 /* 0xbdc0 */;
                12145: data_o = 32'h00000000 /* 0xbdc4 */;
                12146: data_o = 32'h00000000 /* 0xbdc8 */;
                12147: data_o = 32'h00000000 /* 0xbdcc */;
                12148: data_o = 32'h00000000 /* 0xbdd0 */;
                12149: data_o = 32'h00000000 /* 0xbdd4 */;
                12150: data_o = 32'h00000000 /* 0xbdd8 */;
                12151: data_o = 32'h00000000 /* 0xbddc */;
                12152: data_o = 32'h00000000 /* 0xbde0 */;
                12153: data_o = 32'h00000000 /* 0xbde4 */;
                12154: data_o = 32'h00000000 /* 0xbde8 */;
                12155: data_o = 32'h00000000 /* 0xbdec */;
                12156: data_o = 32'h00000000 /* 0xbdf0 */;
                12157: data_o = 32'h00000000 /* 0xbdf4 */;
                12158: data_o = 32'h00000000 /* 0xbdf8 */;
                12159: data_o = 32'h00000000 /* 0xbdfc */;
                12160: data_o = 32'h00000000 /* 0xbe00 */;
                12161: data_o = 32'h00000000 /* 0xbe04 */;
                12162: data_o = 32'h00000000 /* 0xbe08 */;
                12163: data_o = 32'h00000000 /* 0xbe0c */;
                12164: data_o = 32'h00000000 /* 0xbe10 */;
                12165: data_o = 32'h00000000 /* 0xbe14 */;
                12166: data_o = 32'h00000000 /* 0xbe18 */;
                12167: data_o = 32'h00000000 /* 0xbe1c */;
                12168: data_o = 32'h00000000 /* 0xbe20 */;
                12169: data_o = 32'h00000000 /* 0xbe24 */;
                12170: data_o = 32'h00000000 /* 0xbe28 */;
                12171: data_o = 32'h00000000 /* 0xbe2c */;
                12172: data_o = 32'h00000000 /* 0xbe30 */;
                12173: data_o = 32'h00000000 /* 0xbe34 */;
                12174: data_o = 32'h00000000 /* 0xbe38 */;
                12175: data_o = 32'h00000000 /* 0xbe3c */;
                12176: data_o = 32'h00000000 /* 0xbe40 */;
                12177: data_o = 32'h00000000 /* 0xbe44 */;
                12178: data_o = 32'h00000000 /* 0xbe48 */;
                12179: data_o = 32'h00000000 /* 0xbe4c */;
                12180: data_o = 32'h00000000 /* 0xbe50 */;
                12181: data_o = 32'h00000000 /* 0xbe54 */;
                12182: data_o = 32'h00000000 /* 0xbe58 */;
                12183: data_o = 32'h00000000 /* 0xbe5c */;
                12184: data_o = 32'h00000000 /* 0xbe60 */;
                12185: data_o = 32'h00000000 /* 0xbe64 */;
                12186: data_o = 32'h00000000 /* 0xbe68 */;
                12187: data_o = 32'h00000000 /* 0xbe6c */;
                12188: data_o = 32'h00000000 /* 0xbe70 */;
                12189: data_o = 32'h00000000 /* 0xbe74 */;
                12190: data_o = 32'h00000000 /* 0xbe78 */;
                12191: data_o = 32'h00000000 /* 0xbe7c */;
                12192: data_o = 32'h00000000 /* 0xbe80 */;
                12193: data_o = 32'h00000000 /* 0xbe84 */;
                12194: data_o = 32'h00000000 /* 0xbe88 */;
                12195: data_o = 32'h00000000 /* 0xbe8c */;
                12196: data_o = 32'h00000000 /* 0xbe90 */;
                12197: data_o = 32'h00000000 /* 0xbe94 */;
                12198: data_o = 32'h00000000 /* 0xbe98 */;
                12199: data_o = 32'h00000000 /* 0xbe9c */;
                12200: data_o = 32'h00000000 /* 0xbea0 */;
                12201: data_o = 32'h00000000 /* 0xbea4 */;
                12202: data_o = 32'h00000000 /* 0xbea8 */;
                12203: data_o = 32'h00000000 /* 0xbeac */;
                12204: data_o = 32'h00000000 /* 0xbeb0 */;
                12205: data_o = 32'h00000000 /* 0xbeb4 */;
                12206: data_o = 32'h00000000 /* 0xbeb8 */;
                12207: data_o = 32'h00000000 /* 0xbebc */;
                12208: data_o = 32'h00000000 /* 0xbec0 */;
                12209: data_o = 32'h00000000 /* 0xbec4 */;
                12210: data_o = 32'h00000000 /* 0xbec8 */;
                12211: data_o = 32'h00000000 /* 0xbecc */;
                12212: data_o = 32'h00000000 /* 0xbed0 */;
                12213: data_o = 32'h00000000 /* 0xbed4 */;
                12214: data_o = 32'h00000000 /* 0xbed8 */;
                12215: data_o = 32'h00000000 /* 0xbedc */;
                12216: data_o = 32'h00000000 /* 0xbee0 */;
                12217: data_o = 32'h00000000 /* 0xbee4 */;
                12218: data_o = 32'h00000000 /* 0xbee8 */;
                12219: data_o = 32'h00000000 /* 0xbeec */;
                12220: data_o = 32'h00000000 /* 0xbef0 */;
                12221: data_o = 32'h00000000 /* 0xbef4 */;
                12222: data_o = 32'h00000000 /* 0xbef8 */;
                12223: data_o = 32'h00000000 /* 0xbefc */;
                12224: data_o = 32'h00000000 /* 0xbf00 */;
                12225: data_o = 32'h00000000 /* 0xbf04 */;
                12226: data_o = 32'h00000000 /* 0xbf08 */;
                12227: data_o = 32'h00000000 /* 0xbf0c */;
                12228: data_o = 32'h00000000 /* 0xbf10 */;
                12229: data_o = 32'h00000000 /* 0xbf14 */;
                12230: data_o = 32'h00000000 /* 0xbf18 */;
                12231: data_o = 32'h00000000 /* 0xbf1c */;
                12232: data_o = 32'h00000000 /* 0xbf20 */;
                12233: data_o = 32'h00000000 /* 0xbf24 */;
                12234: data_o = 32'h00000000 /* 0xbf28 */;
                12235: data_o = 32'h00000000 /* 0xbf2c */;
                12236: data_o = 32'h00000000 /* 0xbf30 */;
                12237: data_o = 32'h00000000 /* 0xbf34 */;
                12238: data_o = 32'h00000000 /* 0xbf38 */;
                12239: data_o = 32'h00000000 /* 0xbf3c */;
                12240: data_o = 32'h00000000 /* 0xbf40 */;
                12241: data_o = 32'h00000000 /* 0xbf44 */;
                12242: data_o = 32'h00000000 /* 0xbf48 */;
                12243: data_o = 32'h00000000 /* 0xbf4c */;
                12244: data_o = 32'h00000000 /* 0xbf50 */;
                12245: data_o = 32'h00000000 /* 0xbf54 */;
                12246: data_o = 32'h00000000 /* 0xbf58 */;
                12247: data_o = 32'h00000000 /* 0xbf5c */;
                12248: data_o = 32'h00000000 /* 0xbf60 */;
                12249: data_o = 32'h00000000 /* 0xbf64 */;
                12250: data_o = 32'h00000000 /* 0xbf68 */;
                12251: data_o = 32'h00000000 /* 0xbf6c */;
                12252: data_o = 32'h00000000 /* 0xbf70 */;
                12253: data_o = 32'h00000000 /* 0xbf74 */;
                12254: data_o = 32'h00000000 /* 0xbf78 */;
                12255: data_o = 32'h00000000 /* 0xbf7c */;
                12256: data_o = 32'h00000000 /* 0xbf80 */;
                12257: data_o = 32'h00000000 /* 0xbf84 */;
                12258: data_o = 32'h00000000 /* 0xbf88 */;
                12259: data_o = 32'h00000000 /* 0xbf8c */;
                12260: data_o = 32'h00000000 /* 0xbf90 */;
                12261: data_o = 32'h00000000 /* 0xbf94 */;
                12262: data_o = 32'h00000000 /* 0xbf98 */;
                12263: data_o = 32'h00000000 /* 0xbf9c */;
                12264: data_o = 32'h00000000 /* 0xbfa0 */;
                12265: data_o = 32'h00000000 /* 0xbfa4 */;
                12266: data_o = 32'h00000000 /* 0xbfa8 */;
                12267: data_o = 32'h00000000 /* 0xbfac */;
                12268: data_o = 32'h00000000 /* 0xbfb0 */;
                12269: data_o = 32'h00000000 /* 0xbfb4 */;
                12270: data_o = 32'h00000000 /* 0xbfb8 */;
                12271: data_o = 32'h00000000 /* 0xbfbc */;
                12272: data_o = 32'h00000000 /* 0xbfc0 */;
                12273: data_o = 32'h00000000 /* 0xbfc4 */;
                12274: data_o = 32'h00000000 /* 0xbfc8 */;
                12275: data_o = 32'h00000000 /* 0xbfcc */;
                12276: data_o = 32'h00000000 /* 0xbfd0 */;
                12277: data_o = 32'h00000000 /* 0xbfd4 */;
                12278: data_o = 32'h00000000 /* 0xbfd8 */;
                12279: data_o = 32'h00000000 /* 0xbfdc */;
                12280: data_o = 32'h00000000 /* 0xbfe0 */;
                12281: data_o = 32'h00000000 /* 0xbfe4 */;
                12282: data_o = 32'h00000000 /* 0xbfe8 */;
                12283: data_o = 32'h00000000 /* 0xbfec */;
                12284: data_o = 32'h00000000 /* 0xbff0 */;
                12285: data_o = 32'h00000000 /* 0xbff4 */;
                12286: data_o = 32'h00000000 /* 0xbff8 */;
                12287: data_o = 32'h00000000 /* 0xbffc */;
                12288: data_o = 32'h00000000 /* 0xc000 */;
                12289: data_o = 32'h00000000 /* 0xc004 */;
                12290: data_o = 32'h00000000 /* 0xc008 */;
                12291: data_o = 32'h00000000 /* 0xc00c */;
                12292: data_o = 32'h00000000 /* 0xc010 */;
                12293: data_o = 32'h00000000 /* 0xc014 */;
                12294: data_o = 32'h00000000 /* 0xc018 */;
                12295: data_o = 32'h00000000 /* 0xc01c */;
                12296: data_o = 32'h00000000 /* 0xc020 */;
                12297: data_o = 32'h00000000 /* 0xc024 */;
                12298: data_o = 32'h00000000 /* 0xc028 */;
                12299: data_o = 32'h00000000 /* 0xc02c */;
                12300: data_o = 32'h00000000 /* 0xc030 */;
                12301: data_o = 32'h00000000 /* 0xc034 */;
                12302: data_o = 32'h00000000 /* 0xc038 */;
                12303: data_o = 32'h00000000 /* 0xc03c */;
                12304: data_o = 32'h00000000 /* 0xc040 */;
                12305: data_o = 32'h00000000 /* 0xc044 */;
                12306: data_o = 32'h00000000 /* 0xc048 */;
                12307: data_o = 32'h00000000 /* 0xc04c */;
                12308: data_o = 32'h00000000 /* 0xc050 */;
                12309: data_o = 32'h00000000 /* 0xc054 */;
                12310: data_o = 32'h00000000 /* 0xc058 */;
                12311: data_o = 32'h00000000 /* 0xc05c */;
                12312: data_o = 32'h00000000 /* 0xc060 */;
                12313: data_o = 32'h00000000 /* 0xc064 */;
                12314: data_o = 32'h00000000 /* 0xc068 */;
                12315: data_o = 32'h00000000 /* 0xc06c */;
                12316: data_o = 32'h00000000 /* 0xc070 */;
                12317: data_o = 32'h00000000 /* 0xc074 */;
                12318: data_o = 32'h00000000 /* 0xc078 */;
                12319: data_o = 32'h00000000 /* 0xc07c */;
                12320: data_o = 32'h00000000 /* 0xc080 */;
                12321: data_o = 32'h00000000 /* 0xc084 */;
                12322: data_o = 32'h00000000 /* 0xc088 */;
                12323: data_o = 32'h00000000 /* 0xc08c */;
                12324: data_o = 32'h00000000 /* 0xc090 */;
                12325: data_o = 32'h00000000 /* 0xc094 */;
                12326: data_o = 32'h00000000 /* 0xc098 */;
                12327: data_o = 32'h00000000 /* 0xc09c */;
                12328: data_o = 32'h00000000 /* 0xc0a0 */;
                12329: data_o = 32'h00000000 /* 0xc0a4 */;
                12330: data_o = 32'h00000000 /* 0xc0a8 */;
                12331: data_o = 32'h00000000 /* 0xc0ac */;
                12332: data_o = 32'h00000000 /* 0xc0b0 */;
                12333: data_o = 32'h00000000 /* 0xc0b4 */;
                12334: data_o = 32'h00000000 /* 0xc0b8 */;
                12335: data_o = 32'h00000000 /* 0xc0bc */;
                12336: data_o = 32'h00000000 /* 0xc0c0 */;
                12337: data_o = 32'h00000000 /* 0xc0c4 */;
                12338: data_o = 32'h00000000 /* 0xc0c8 */;
                12339: data_o = 32'h00000000 /* 0xc0cc */;
                12340: data_o = 32'h00000000 /* 0xc0d0 */;
                12341: data_o = 32'h00000000 /* 0xc0d4 */;
                12342: data_o = 32'h00000000 /* 0xc0d8 */;
                12343: data_o = 32'h00000000 /* 0xc0dc */;
                12344: data_o = 32'h00000000 /* 0xc0e0 */;
                12345: data_o = 32'h00000000 /* 0xc0e4 */;
                12346: data_o = 32'h00000000 /* 0xc0e8 */;
                12347: data_o = 32'h00000000 /* 0xc0ec */;
                12348: data_o = 32'h00000000 /* 0xc0f0 */;
                12349: data_o = 32'h00000000 /* 0xc0f4 */;
                12350: data_o = 32'h00000000 /* 0xc0f8 */;
                12351: data_o = 32'h00000000 /* 0xc0fc */;
                12352: data_o = 32'h00000000 /* 0xc100 */;
                12353: data_o = 32'h00000000 /* 0xc104 */;
                12354: data_o = 32'h00000000 /* 0xc108 */;
                12355: data_o = 32'h00000000 /* 0xc10c */;
                12356: data_o = 32'h00000000 /* 0xc110 */;
                12357: data_o = 32'h00000000 /* 0xc114 */;
                12358: data_o = 32'h00000000 /* 0xc118 */;
                12359: data_o = 32'h00000000 /* 0xc11c */;
                12360: data_o = 32'h00000000 /* 0xc120 */;
                12361: data_o = 32'h00000000 /* 0xc124 */;
                12362: data_o = 32'h00000000 /* 0xc128 */;
                12363: data_o = 32'h00000000 /* 0xc12c */;
                12364: data_o = 32'h00000000 /* 0xc130 */;
                12365: data_o = 32'h00000000 /* 0xc134 */;
                12366: data_o = 32'h00000000 /* 0xc138 */;
                12367: data_o = 32'h00000000 /* 0xc13c */;
                12368: data_o = 32'h00000000 /* 0xc140 */;
                12369: data_o = 32'h00000000 /* 0xc144 */;
                12370: data_o = 32'h00000000 /* 0xc148 */;
                12371: data_o = 32'h00000000 /* 0xc14c */;
                12372: data_o = 32'h00000000 /* 0xc150 */;
                12373: data_o = 32'h00000000 /* 0xc154 */;
                12374: data_o = 32'h00000000 /* 0xc158 */;
                12375: data_o = 32'h00000000 /* 0xc15c */;
                12376: data_o = 32'h00000000 /* 0xc160 */;
                12377: data_o = 32'h00000000 /* 0xc164 */;
                12378: data_o = 32'h00000000 /* 0xc168 */;
                12379: data_o = 32'h00000000 /* 0xc16c */;
                12380: data_o = 32'h00000000 /* 0xc170 */;
                12381: data_o = 32'h00000000 /* 0xc174 */;
                12382: data_o = 32'h00000000 /* 0xc178 */;
                12383: data_o = 32'h00000000 /* 0xc17c */;
                12384: data_o = 32'h00000000 /* 0xc180 */;
                12385: data_o = 32'h00000000 /* 0xc184 */;
                12386: data_o = 32'h00000000 /* 0xc188 */;
                12387: data_o = 32'h00000000 /* 0xc18c */;
                12388: data_o = 32'h00000000 /* 0xc190 */;
                12389: data_o = 32'h00000000 /* 0xc194 */;
                12390: data_o = 32'h00000000 /* 0xc198 */;
                12391: data_o = 32'h00000000 /* 0xc19c */;
                12392: data_o = 32'h00000000 /* 0xc1a0 */;
                12393: data_o = 32'h00000000 /* 0xc1a4 */;
                12394: data_o = 32'h00000000 /* 0xc1a8 */;
                12395: data_o = 32'h00000000 /* 0xc1ac */;
                12396: data_o = 32'h00000000 /* 0xc1b0 */;
                12397: data_o = 32'h00000000 /* 0xc1b4 */;
                12398: data_o = 32'h00000000 /* 0xc1b8 */;
                12399: data_o = 32'h00000000 /* 0xc1bc */;
                12400: data_o = 32'h00000000 /* 0xc1c0 */;
                12401: data_o = 32'h00000000 /* 0xc1c4 */;
                12402: data_o = 32'h00000000 /* 0xc1c8 */;
                12403: data_o = 32'h00000000 /* 0xc1cc */;
                12404: data_o = 32'h00000000 /* 0xc1d0 */;
                12405: data_o = 32'h00000000 /* 0xc1d4 */;
                12406: data_o = 32'h00000000 /* 0xc1d8 */;
                12407: data_o = 32'h00000000 /* 0xc1dc */;
                12408: data_o = 32'h00000000 /* 0xc1e0 */;
                12409: data_o = 32'h00000000 /* 0xc1e4 */;
                12410: data_o = 32'h00000000 /* 0xc1e8 */;
                12411: data_o = 32'h00000000 /* 0xc1ec */;
                12412: data_o = 32'h00000000 /* 0xc1f0 */;
                12413: data_o = 32'h00000000 /* 0xc1f4 */;
                12414: data_o = 32'h00000000 /* 0xc1f8 */;
                12415: data_o = 32'h00000000 /* 0xc1fc */;
                12416: data_o = 32'h00000000 /* 0xc200 */;
                12417: data_o = 32'h00000000 /* 0xc204 */;
                12418: data_o = 32'h00000000 /* 0xc208 */;
                12419: data_o = 32'h00000000 /* 0xc20c */;
                12420: data_o = 32'h00000000 /* 0xc210 */;
                12421: data_o = 32'h00000000 /* 0xc214 */;
                12422: data_o = 32'h00000000 /* 0xc218 */;
                12423: data_o = 32'h00000000 /* 0xc21c */;
                12424: data_o = 32'h00000000 /* 0xc220 */;
                12425: data_o = 32'h00000000 /* 0xc224 */;
                12426: data_o = 32'h00000000 /* 0xc228 */;
                12427: data_o = 32'h00000000 /* 0xc22c */;
                12428: data_o = 32'h00000000 /* 0xc230 */;
                12429: data_o = 32'h00000000 /* 0xc234 */;
                12430: data_o = 32'h00000000 /* 0xc238 */;
                12431: data_o = 32'h00000000 /* 0xc23c */;
                12432: data_o = 32'h00000000 /* 0xc240 */;
                12433: data_o = 32'h00000000 /* 0xc244 */;
                12434: data_o = 32'h00000000 /* 0xc248 */;
                12435: data_o = 32'h00000000 /* 0xc24c */;
                12436: data_o = 32'h00000000 /* 0xc250 */;
                12437: data_o = 32'h00000000 /* 0xc254 */;
                12438: data_o = 32'h00000000 /* 0xc258 */;
                12439: data_o = 32'h00000000 /* 0xc25c */;
                12440: data_o = 32'h00000000 /* 0xc260 */;
                12441: data_o = 32'h00000000 /* 0xc264 */;
                12442: data_o = 32'h00000000 /* 0xc268 */;
                12443: data_o = 32'h00000000 /* 0xc26c */;
                12444: data_o = 32'h00000000 /* 0xc270 */;
                12445: data_o = 32'h00000000 /* 0xc274 */;
                12446: data_o = 32'h00000000 /* 0xc278 */;
                12447: data_o = 32'h00000000 /* 0xc27c */;
                12448: data_o = 32'h00000000 /* 0xc280 */;
                12449: data_o = 32'h00000000 /* 0xc284 */;
                12450: data_o = 32'h00000000 /* 0xc288 */;
                12451: data_o = 32'h00000000 /* 0xc28c */;
                12452: data_o = 32'h00000000 /* 0xc290 */;
                12453: data_o = 32'h00000000 /* 0xc294 */;
                12454: data_o = 32'h00000000 /* 0xc298 */;
                12455: data_o = 32'h00000000 /* 0xc29c */;
                12456: data_o = 32'h00000000 /* 0xc2a0 */;
                12457: data_o = 32'h00000000 /* 0xc2a4 */;
                12458: data_o = 32'h00000000 /* 0xc2a8 */;
                12459: data_o = 32'h00000000 /* 0xc2ac */;
                12460: data_o = 32'h00000000 /* 0xc2b0 */;
                12461: data_o = 32'h00000000 /* 0xc2b4 */;
                12462: data_o = 32'h00000000 /* 0xc2b8 */;
                12463: data_o = 32'h00000000 /* 0xc2bc */;
                12464: data_o = 32'h00000000 /* 0xc2c0 */;
                12465: data_o = 32'h00000000 /* 0xc2c4 */;
                12466: data_o = 32'h00000000 /* 0xc2c8 */;
                12467: data_o = 32'h00000000 /* 0xc2cc */;
                12468: data_o = 32'h00000000 /* 0xc2d0 */;
                12469: data_o = 32'h00000000 /* 0xc2d4 */;
                12470: data_o = 32'h00000000 /* 0xc2d8 */;
                12471: data_o = 32'h00000000 /* 0xc2dc */;
                12472: data_o = 32'h00000000 /* 0xc2e0 */;
                12473: data_o = 32'h00000000 /* 0xc2e4 */;
                12474: data_o = 32'h00000000 /* 0xc2e8 */;
                12475: data_o = 32'h00000000 /* 0xc2ec */;
                12476: data_o = 32'h00000000 /* 0xc2f0 */;
                12477: data_o = 32'h00000000 /* 0xc2f4 */;
                12478: data_o = 32'h00000000 /* 0xc2f8 */;
                12479: data_o = 32'h00000000 /* 0xc2fc */;
                12480: data_o = 32'h00000000 /* 0xc300 */;
                12481: data_o = 32'h00000000 /* 0xc304 */;
                12482: data_o = 32'h00000000 /* 0xc308 */;
                12483: data_o = 32'h00000000 /* 0xc30c */;
                12484: data_o = 32'h00000000 /* 0xc310 */;
                12485: data_o = 32'h00000000 /* 0xc314 */;
                12486: data_o = 32'h00000000 /* 0xc318 */;
                12487: data_o = 32'h00000000 /* 0xc31c */;
                12488: data_o = 32'h00000000 /* 0xc320 */;
                12489: data_o = 32'h00000000 /* 0xc324 */;
                12490: data_o = 32'h00000000 /* 0xc328 */;
                12491: data_o = 32'h00000000 /* 0xc32c */;
                12492: data_o = 32'h00000000 /* 0xc330 */;
                12493: data_o = 32'h00000000 /* 0xc334 */;
                12494: data_o = 32'h00000000 /* 0xc338 */;
                12495: data_o = 32'h00000000 /* 0xc33c */;
                12496: data_o = 32'h00000000 /* 0xc340 */;
                12497: data_o = 32'h00000000 /* 0xc344 */;
                12498: data_o = 32'h00000000 /* 0xc348 */;
                12499: data_o = 32'h00000000 /* 0xc34c */;
                12500: data_o = 32'h00000000 /* 0xc350 */;
                12501: data_o = 32'h00000000 /* 0xc354 */;
                12502: data_o = 32'h00000000 /* 0xc358 */;
                12503: data_o = 32'h00000000 /* 0xc35c */;
                12504: data_o = 32'h00000000 /* 0xc360 */;
                12505: data_o = 32'h00000000 /* 0xc364 */;
                12506: data_o = 32'h00000000 /* 0xc368 */;
                12507: data_o = 32'h00000000 /* 0xc36c */;
                12508: data_o = 32'h00000000 /* 0xc370 */;
                12509: data_o = 32'h00000000 /* 0xc374 */;
                12510: data_o = 32'h00000000 /* 0xc378 */;
                12511: data_o = 32'h00000000 /* 0xc37c */;
                12512: data_o = 32'h00000000 /* 0xc380 */;
                12513: data_o = 32'h00000000 /* 0xc384 */;
                12514: data_o = 32'h00000000 /* 0xc388 */;
                12515: data_o = 32'h00000000 /* 0xc38c */;
                12516: data_o = 32'h00000000 /* 0xc390 */;
                12517: data_o = 32'h00000000 /* 0xc394 */;
                12518: data_o = 32'h00000000 /* 0xc398 */;
                12519: data_o = 32'h00000000 /* 0xc39c */;
                12520: data_o = 32'h00000000 /* 0xc3a0 */;
                12521: data_o = 32'h00000000 /* 0xc3a4 */;
                12522: data_o = 32'h00000000 /* 0xc3a8 */;
                12523: data_o = 32'h00000000 /* 0xc3ac */;
                12524: data_o = 32'h00000000 /* 0xc3b0 */;
                12525: data_o = 32'h00000000 /* 0xc3b4 */;
                12526: data_o = 32'h00000000 /* 0xc3b8 */;
                12527: data_o = 32'h00000000 /* 0xc3bc */;
                12528: data_o = 32'h00000000 /* 0xc3c0 */;
                12529: data_o = 32'h00000000 /* 0xc3c4 */;
                12530: data_o = 32'h00000000 /* 0xc3c8 */;
                12531: data_o = 32'h00000000 /* 0xc3cc */;
                12532: data_o = 32'h00000000 /* 0xc3d0 */;
                12533: data_o = 32'h00000000 /* 0xc3d4 */;
                12534: data_o = 32'h00000000 /* 0xc3d8 */;
                12535: data_o = 32'h00000000 /* 0xc3dc */;
                12536: data_o = 32'h00000000 /* 0xc3e0 */;
                12537: data_o = 32'h00000000 /* 0xc3e4 */;
                12538: data_o = 32'h00000000 /* 0xc3e8 */;
                12539: data_o = 32'h00000000 /* 0xc3ec */;
                12540: data_o = 32'h00000000 /* 0xc3f0 */;
                12541: data_o = 32'h00000000 /* 0xc3f4 */;
                12542: data_o = 32'h00000000 /* 0xc3f8 */;
                12543: data_o = 32'h00000000 /* 0xc3fc */;
                12544: data_o = 32'h00000000 /* 0xc400 */;
                12545: data_o = 32'h00000000 /* 0xc404 */;
                12546: data_o = 32'h00000000 /* 0xc408 */;
                12547: data_o = 32'h00000000 /* 0xc40c */;
                12548: data_o = 32'h00000000 /* 0xc410 */;
                12549: data_o = 32'h00000000 /* 0xc414 */;
                12550: data_o = 32'h00000000 /* 0xc418 */;
                12551: data_o = 32'h00000000 /* 0xc41c */;
                12552: data_o = 32'h00000000 /* 0xc420 */;
                12553: data_o = 32'h00000000 /* 0xc424 */;
                12554: data_o = 32'h00000000 /* 0xc428 */;
                12555: data_o = 32'h00000000 /* 0xc42c */;
                12556: data_o = 32'h00000000 /* 0xc430 */;
                12557: data_o = 32'h00000000 /* 0xc434 */;
                12558: data_o = 32'h00000000 /* 0xc438 */;
                12559: data_o = 32'h00000000 /* 0xc43c */;
                12560: data_o = 32'h00000000 /* 0xc440 */;
                12561: data_o = 32'h00000000 /* 0xc444 */;
                12562: data_o = 32'h00000000 /* 0xc448 */;
                12563: data_o = 32'h00000000 /* 0xc44c */;
                12564: data_o = 32'h00000000 /* 0xc450 */;
                12565: data_o = 32'h00000000 /* 0xc454 */;
                12566: data_o = 32'h00000000 /* 0xc458 */;
                12567: data_o = 32'h00000000 /* 0xc45c */;
                12568: data_o = 32'h00000000 /* 0xc460 */;
                12569: data_o = 32'h00000000 /* 0xc464 */;
                12570: data_o = 32'h00000000 /* 0xc468 */;
                12571: data_o = 32'h00000000 /* 0xc46c */;
                12572: data_o = 32'h00000000 /* 0xc470 */;
                12573: data_o = 32'h00000000 /* 0xc474 */;
                12574: data_o = 32'h00000000 /* 0xc478 */;
                12575: data_o = 32'h00000000 /* 0xc47c */;
                12576: data_o = 32'h00000000 /* 0xc480 */;
                12577: data_o = 32'h00000000 /* 0xc484 */;
                12578: data_o = 32'h00000000 /* 0xc488 */;
                12579: data_o = 32'h00000000 /* 0xc48c */;
                12580: data_o = 32'h00000000 /* 0xc490 */;
                12581: data_o = 32'h00000000 /* 0xc494 */;
                12582: data_o = 32'h00000000 /* 0xc498 */;
                12583: data_o = 32'h00000000 /* 0xc49c */;
                12584: data_o = 32'h00000000 /* 0xc4a0 */;
                12585: data_o = 32'h00000000 /* 0xc4a4 */;
                12586: data_o = 32'h00000000 /* 0xc4a8 */;
                12587: data_o = 32'h00000000 /* 0xc4ac */;
                12588: data_o = 32'h00000000 /* 0xc4b0 */;
                12589: data_o = 32'h00000000 /* 0xc4b4 */;
                12590: data_o = 32'h00000000 /* 0xc4b8 */;
                12591: data_o = 32'h00000000 /* 0xc4bc */;
                12592: data_o = 32'h00000000 /* 0xc4c0 */;
                12593: data_o = 32'h00000000 /* 0xc4c4 */;
                12594: data_o = 32'h00000000 /* 0xc4c8 */;
                12595: data_o = 32'h00000000 /* 0xc4cc */;
                12596: data_o = 32'h00000000 /* 0xc4d0 */;
                12597: data_o = 32'h00000000 /* 0xc4d4 */;
                12598: data_o = 32'h00000000 /* 0xc4d8 */;
                12599: data_o = 32'h00000000 /* 0xc4dc */;
                12600: data_o = 32'h00000000 /* 0xc4e0 */;
                12601: data_o = 32'h00000000 /* 0xc4e4 */;
                12602: data_o = 32'h00000000 /* 0xc4e8 */;
                12603: data_o = 32'h00000000 /* 0xc4ec */;
                12604: data_o = 32'h00000000 /* 0xc4f0 */;
                12605: data_o = 32'h00000000 /* 0xc4f4 */;
                12606: data_o = 32'h00000000 /* 0xc4f8 */;
                12607: data_o = 32'h00000000 /* 0xc4fc */;
                12608: data_o = 32'h00000000 /* 0xc500 */;
                12609: data_o = 32'h00000000 /* 0xc504 */;
                12610: data_o = 32'h00000000 /* 0xc508 */;
                12611: data_o = 32'h00000000 /* 0xc50c */;
                12612: data_o = 32'h00000000 /* 0xc510 */;
                12613: data_o = 32'h00000000 /* 0xc514 */;
                12614: data_o = 32'h00000000 /* 0xc518 */;
                12615: data_o = 32'h00000000 /* 0xc51c */;
                12616: data_o = 32'h00000000 /* 0xc520 */;
                12617: data_o = 32'h00000000 /* 0xc524 */;
                12618: data_o = 32'h00000000 /* 0xc528 */;
                12619: data_o = 32'h00000000 /* 0xc52c */;
                12620: data_o = 32'h00000000 /* 0xc530 */;
                12621: data_o = 32'h00000000 /* 0xc534 */;
                12622: data_o = 32'h00000000 /* 0xc538 */;
                12623: data_o = 32'h00000000 /* 0xc53c */;
                12624: data_o = 32'h00000000 /* 0xc540 */;
                12625: data_o = 32'h00000000 /* 0xc544 */;
                12626: data_o = 32'h00000000 /* 0xc548 */;
                12627: data_o = 32'h00000000 /* 0xc54c */;
                12628: data_o = 32'h00000000 /* 0xc550 */;
                12629: data_o = 32'h00000000 /* 0xc554 */;
                12630: data_o = 32'h00000000 /* 0xc558 */;
                12631: data_o = 32'h00000000 /* 0xc55c */;
                12632: data_o = 32'h00000000 /* 0xc560 */;
                12633: data_o = 32'h00000000 /* 0xc564 */;
                12634: data_o = 32'h00000000 /* 0xc568 */;
                12635: data_o = 32'h00000000 /* 0xc56c */;
                12636: data_o = 32'h00000000 /* 0xc570 */;
                12637: data_o = 32'h00000000 /* 0xc574 */;
                12638: data_o = 32'h00000000 /* 0xc578 */;
                12639: data_o = 32'h00000000 /* 0xc57c */;
                12640: data_o = 32'h00000000 /* 0xc580 */;
                12641: data_o = 32'h00000000 /* 0xc584 */;
                12642: data_o = 32'h00000000 /* 0xc588 */;
                12643: data_o = 32'h00000000 /* 0xc58c */;
                12644: data_o = 32'h00000000 /* 0xc590 */;
                12645: data_o = 32'h00000000 /* 0xc594 */;
                12646: data_o = 32'h00000000 /* 0xc598 */;
                12647: data_o = 32'h00000000 /* 0xc59c */;
                12648: data_o = 32'h00000000 /* 0xc5a0 */;
                12649: data_o = 32'h00000000 /* 0xc5a4 */;
                12650: data_o = 32'h00000000 /* 0xc5a8 */;
                12651: data_o = 32'h00000000 /* 0xc5ac */;
                12652: data_o = 32'h00000000 /* 0xc5b0 */;
                12653: data_o = 32'h00000000 /* 0xc5b4 */;
                12654: data_o = 32'h00000000 /* 0xc5b8 */;
                12655: data_o = 32'h00000000 /* 0xc5bc */;
                12656: data_o = 32'h00000000 /* 0xc5c0 */;
                12657: data_o = 32'h00000000 /* 0xc5c4 */;
                12658: data_o = 32'h00000000 /* 0xc5c8 */;
                12659: data_o = 32'h00000000 /* 0xc5cc */;
                12660: data_o = 32'h00000000 /* 0xc5d0 */;
                12661: data_o = 32'h00000000 /* 0xc5d4 */;
                12662: data_o = 32'h00000000 /* 0xc5d8 */;
                12663: data_o = 32'h00000000 /* 0xc5dc */;
                12664: data_o = 32'h00000000 /* 0xc5e0 */;
                12665: data_o = 32'h00000000 /* 0xc5e4 */;
                12666: data_o = 32'h00000000 /* 0xc5e8 */;
                12667: data_o = 32'h00000000 /* 0xc5ec */;
                12668: data_o = 32'h00000000 /* 0xc5f0 */;
                12669: data_o = 32'h00000000 /* 0xc5f4 */;
                12670: data_o = 32'h00000000 /* 0xc5f8 */;
                12671: data_o = 32'h00000000 /* 0xc5fc */;
                12672: data_o = 32'h00000000 /* 0xc600 */;
                12673: data_o = 32'h00000000 /* 0xc604 */;
                12674: data_o = 32'h00000000 /* 0xc608 */;
                12675: data_o = 32'h00000000 /* 0xc60c */;
                12676: data_o = 32'h00000000 /* 0xc610 */;
                12677: data_o = 32'h00000000 /* 0xc614 */;
                12678: data_o = 32'h00000000 /* 0xc618 */;
                12679: data_o = 32'h00000000 /* 0xc61c */;
                12680: data_o = 32'h00000000 /* 0xc620 */;
                12681: data_o = 32'h00000000 /* 0xc624 */;
                12682: data_o = 32'h00000000 /* 0xc628 */;
                12683: data_o = 32'h00000000 /* 0xc62c */;
                12684: data_o = 32'h00000000 /* 0xc630 */;
                12685: data_o = 32'h00000000 /* 0xc634 */;
                12686: data_o = 32'h00000000 /* 0xc638 */;
                12687: data_o = 32'h00000000 /* 0xc63c */;
                12688: data_o = 32'h00000000 /* 0xc640 */;
                12689: data_o = 32'h00000000 /* 0xc644 */;
                12690: data_o = 32'h00000000 /* 0xc648 */;
                12691: data_o = 32'h00000000 /* 0xc64c */;
                12692: data_o = 32'h00000000 /* 0xc650 */;
                12693: data_o = 32'h00000000 /* 0xc654 */;
                12694: data_o = 32'h00000000 /* 0xc658 */;
                12695: data_o = 32'h00000000 /* 0xc65c */;
                12696: data_o = 32'h00000000 /* 0xc660 */;
                12697: data_o = 32'h00000000 /* 0xc664 */;
                12698: data_o = 32'h00000000 /* 0xc668 */;
                12699: data_o = 32'h00000000 /* 0xc66c */;
                12700: data_o = 32'h00000000 /* 0xc670 */;
                12701: data_o = 32'h00000000 /* 0xc674 */;
                12702: data_o = 32'h00000000 /* 0xc678 */;
                12703: data_o = 32'h00000000 /* 0xc67c */;
                12704: data_o = 32'h00000000 /* 0xc680 */;
                12705: data_o = 32'h00000000 /* 0xc684 */;
                12706: data_o = 32'h00000000 /* 0xc688 */;
                12707: data_o = 32'h00000000 /* 0xc68c */;
                12708: data_o = 32'h00000000 /* 0xc690 */;
                12709: data_o = 32'h00000000 /* 0xc694 */;
                12710: data_o = 32'h00000000 /* 0xc698 */;
                12711: data_o = 32'h00000000 /* 0xc69c */;
                12712: data_o = 32'h00000000 /* 0xc6a0 */;
                12713: data_o = 32'h00000000 /* 0xc6a4 */;
                12714: data_o = 32'h00000000 /* 0xc6a8 */;
                12715: data_o = 32'h00000000 /* 0xc6ac */;
                12716: data_o = 32'h00000000 /* 0xc6b0 */;
                12717: data_o = 32'h00000000 /* 0xc6b4 */;
                12718: data_o = 32'h00000000 /* 0xc6b8 */;
                12719: data_o = 32'h00000000 /* 0xc6bc */;
                12720: data_o = 32'h00000000 /* 0xc6c0 */;
                12721: data_o = 32'h00000000 /* 0xc6c4 */;
                12722: data_o = 32'h00000000 /* 0xc6c8 */;
                12723: data_o = 32'h00000000 /* 0xc6cc */;
                12724: data_o = 32'h00000000 /* 0xc6d0 */;
                12725: data_o = 32'h00000000 /* 0xc6d4 */;
                12726: data_o = 32'h00000000 /* 0xc6d8 */;
                12727: data_o = 32'h00000000 /* 0xc6dc */;
                12728: data_o = 32'h00000000 /* 0xc6e0 */;
                12729: data_o = 32'h00000000 /* 0xc6e4 */;
                12730: data_o = 32'h00000000 /* 0xc6e8 */;
                12731: data_o = 32'h00000000 /* 0xc6ec */;
                12732: data_o = 32'h00000000 /* 0xc6f0 */;
                12733: data_o = 32'h00000000 /* 0xc6f4 */;
                12734: data_o = 32'h00000000 /* 0xc6f8 */;
                12735: data_o = 32'h00000000 /* 0xc6fc */;
                12736: data_o = 32'h00000000 /* 0xc700 */;
                12737: data_o = 32'h00000000 /* 0xc704 */;
                12738: data_o = 32'h00000000 /* 0xc708 */;
                12739: data_o = 32'h00000000 /* 0xc70c */;
                12740: data_o = 32'h00000000 /* 0xc710 */;
                12741: data_o = 32'h00000000 /* 0xc714 */;
                12742: data_o = 32'h00000000 /* 0xc718 */;
                12743: data_o = 32'h00000000 /* 0xc71c */;
                12744: data_o = 32'h00000000 /* 0xc720 */;
                12745: data_o = 32'h00000000 /* 0xc724 */;
                12746: data_o = 32'h00000000 /* 0xc728 */;
                12747: data_o = 32'h00000000 /* 0xc72c */;
                12748: data_o = 32'h00000000 /* 0xc730 */;
                12749: data_o = 32'h00000000 /* 0xc734 */;
                12750: data_o = 32'h00000000 /* 0xc738 */;
                12751: data_o = 32'h00000000 /* 0xc73c */;
                12752: data_o = 32'h00000000 /* 0xc740 */;
                12753: data_o = 32'h00000000 /* 0xc744 */;
                12754: data_o = 32'h00000000 /* 0xc748 */;
                12755: data_o = 32'h00000000 /* 0xc74c */;
                12756: data_o = 32'h00000000 /* 0xc750 */;
                12757: data_o = 32'h00000000 /* 0xc754 */;
                12758: data_o = 32'h00000000 /* 0xc758 */;
                12759: data_o = 32'h00000000 /* 0xc75c */;
                12760: data_o = 32'h00000000 /* 0xc760 */;
                12761: data_o = 32'h00000000 /* 0xc764 */;
                12762: data_o = 32'h00000000 /* 0xc768 */;
                12763: data_o = 32'h00000000 /* 0xc76c */;
                12764: data_o = 32'h00000000 /* 0xc770 */;
                12765: data_o = 32'h00000000 /* 0xc774 */;
                12766: data_o = 32'h00000000 /* 0xc778 */;
                12767: data_o = 32'h00000000 /* 0xc77c */;
                12768: data_o = 32'h00000000 /* 0xc780 */;
                12769: data_o = 32'h00000000 /* 0xc784 */;
                12770: data_o = 32'h00000000 /* 0xc788 */;
                12771: data_o = 32'h00000000 /* 0xc78c */;
                12772: data_o = 32'h00000000 /* 0xc790 */;
                12773: data_o = 32'h00000000 /* 0xc794 */;
                12774: data_o = 32'h00000000 /* 0xc798 */;
                12775: data_o = 32'h00000000 /* 0xc79c */;
                12776: data_o = 32'h00000000 /* 0xc7a0 */;
                12777: data_o = 32'h00000000 /* 0xc7a4 */;
                12778: data_o = 32'h00000000 /* 0xc7a8 */;
                12779: data_o = 32'h00000000 /* 0xc7ac */;
                12780: data_o = 32'h00000000 /* 0xc7b0 */;
                12781: data_o = 32'h00000000 /* 0xc7b4 */;
                12782: data_o = 32'h00000000 /* 0xc7b8 */;
                12783: data_o = 32'h00000000 /* 0xc7bc */;
                12784: data_o = 32'h00000000 /* 0xc7c0 */;
                12785: data_o = 32'h00000000 /* 0xc7c4 */;
                12786: data_o = 32'h00000000 /* 0xc7c8 */;
                12787: data_o = 32'h00000000 /* 0xc7cc */;
                12788: data_o = 32'h00000000 /* 0xc7d0 */;
                12789: data_o = 32'h00000000 /* 0xc7d4 */;
                12790: data_o = 32'h00000000 /* 0xc7d8 */;
                12791: data_o = 32'h00000000 /* 0xc7dc */;
                12792: data_o = 32'h00000000 /* 0xc7e0 */;
                12793: data_o = 32'h00000000 /* 0xc7e4 */;
                12794: data_o = 32'h00000000 /* 0xc7e8 */;
                12795: data_o = 32'h00000000 /* 0xc7ec */;
                12796: data_o = 32'h00000000 /* 0xc7f0 */;
                12797: data_o = 32'h00000000 /* 0xc7f4 */;
                12798: data_o = 32'h00000000 /* 0xc7f8 */;
                12799: data_o = 32'h00000000 /* 0xc7fc */;
                12800: data_o = 32'h00000000 /* 0xc800 */;
                12801: data_o = 32'h00000000 /* 0xc804 */;
                12802: data_o = 32'h00000000 /* 0xc808 */;
                12803: data_o = 32'h00000000 /* 0xc80c */;
                12804: data_o = 32'h00000000 /* 0xc810 */;
                12805: data_o = 32'h00000000 /* 0xc814 */;
                12806: data_o = 32'h00000000 /* 0xc818 */;
                12807: data_o = 32'h00000000 /* 0xc81c */;
                12808: data_o = 32'h00000000 /* 0xc820 */;
                12809: data_o = 32'h00000000 /* 0xc824 */;
                12810: data_o = 32'h00000000 /* 0xc828 */;
                12811: data_o = 32'h00000000 /* 0xc82c */;
                12812: data_o = 32'h00000000 /* 0xc830 */;
                12813: data_o = 32'h00000000 /* 0xc834 */;
                12814: data_o = 32'h00000000 /* 0xc838 */;
                12815: data_o = 32'h00000000 /* 0xc83c */;
                12816: data_o = 32'h00000000 /* 0xc840 */;
                12817: data_o = 32'h00000000 /* 0xc844 */;
                12818: data_o = 32'h00000000 /* 0xc848 */;
                12819: data_o = 32'h00000000 /* 0xc84c */;
                12820: data_o = 32'h00000000 /* 0xc850 */;
                12821: data_o = 32'h00000000 /* 0xc854 */;
                12822: data_o = 32'h00000000 /* 0xc858 */;
                12823: data_o = 32'h00000000 /* 0xc85c */;
                12824: data_o = 32'h00000000 /* 0xc860 */;
                12825: data_o = 32'h00000000 /* 0xc864 */;
                12826: data_o = 32'h00000000 /* 0xc868 */;
                12827: data_o = 32'h00000000 /* 0xc86c */;
                12828: data_o = 32'h00000000 /* 0xc870 */;
                12829: data_o = 32'h00000000 /* 0xc874 */;
                12830: data_o = 32'h00000000 /* 0xc878 */;
                12831: data_o = 32'h00000000 /* 0xc87c */;
                12832: data_o = 32'h00000000 /* 0xc880 */;
                12833: data_o = 32'h00000000 /* 0xc884 */;
                12834: data_o = 32'h00000000 /* 0xc888 */;
                12835: data_o = 32'h00000000 /* 0xc88c */;
                12836: data_o = 32'h00000000 /* 0xc890 */;
                12837: data_o = 32'h00000000 /* 0xc894 */;
                12838: data_o = 32'h00000000 /* 0xc898 */;
                12839: data_o = 32'h00000000 /* 0xc89c */;
                12840: data_o = 32'h00000000 /* 0xc8a0 */;
                12841: data_o = 32'h00000000 /* 0xc8a4 */;
                12842: data_o = 32'h00000000 /* 0xc8a8 */;
                12843: data_o = 32'h00000000 /* 0xc8ac */;
                12844: data_o = 32'h00000000 /* 0xc8b0 */;
                12845: data_o = 32'h00000000 /* 0xc8b4 */;
                12846: data_o = 32'h00000000 /* 0xc8b8 */;
                12847: data_o = 32'h00000000 /* 0xc8bc */;
                12848: data_o = 32'h00000000 /* 0xc8c0 */;
                12849: data_o = 32'h00000000 /* 0xc8c4 */;
                12850: data_o = 32'h00000000 /* 0xc8c8 */;
                12851: data_o = 32'h00000000 /* 0xc8cc */;
                12852: data_o = 32'h00000000 /* 0xc8d0 */;
                12853: data_o = 32'h00000000 /* 0xc8d4 */;
                12854: data_o = 32'h00000000 /* 0xc8d8 */;
                12855: data_o = 32'h00000000 /* 0xc8dc */;
                12856: data_o = 32'h00000000 /* 0xc8e0 */;
                12857: data_o = 32'h00000000 /* 0xc8e4 */;
                12858: data_o = 32'h00000000 /* 0xc8e8 */;
                12859: data_o = 32'h00000000 /* 0xc8ec */;
                12860: data_o = 32'h00000000 /* 0xc8f0 */;
                12861: data_o = 32'h00000000 /* 0xc8f4 */;
                12862: data_o = 32'h00000000 /* 0xc8f8 */;
                12863: data_o = 32'h00000000 /* 0xc8fc */;
                12864: data_o = 32'h00000000 /* 0xc900 */;
                12865: data_o = 32'h00000000 /* 0xc904 */;
                12866: data_o = 32'h00000000 /* 0xc908 */;
                12867: data_o = 32'h00000000 /* 0xc90c */;
                12868: data_o = 32'h00000000 /* 0xc910 */;
                12869: data_o = 32'h00000000 /* 0xc914 */;
                12870: data_o = 32'h00000000 /* 0xc918 */;
                12871: data_o = 32'h00000000 /* 0xc91c */;
                12872: data_o = 32'h00000000 /* 0xc920 */;
                12873: data_o = 32'h00000000 /* 0xc924 */;
                12874: data_o = 32'h00000000 /* 0xc928 */;
                12875: data_o = 32'h00000000 /* 0xc92c */;
                12876: data_o = 32'h00000000 /* 0xc930 */;
                12877: data_o = 32'h00000000 /* 0xc934 */;
                12878: data_o = 32'h00000000 /* 0xc938 */;
                12879: data_o = 32'h00000000 /* 0xc93c */;
                12880: data_o = 32'h00000000 /* 0xc940 */;
                12881: data_o = 32'h00000000 /* 0xc944 */;
                12882: data_o = 32'h00000000 /* 0xc948 */;
                12883: data_o = 32'h00000000 /* 0xc94c */;
                12884: data_o = 32'h00000000 /* 0xc950 */;
                12885: data_o = 32'h00000000 /* 0xc954 */;
                12886: data_o = 32'h00000000 /* 0xc958 */;
                12887: data_o = 32'h00000000 /* 0xc95c */;
                12888: data_o = 32'h00000000 /* 0xc960 */;
                12889: data_o = 32'h00000000 /* 0xc964 */;
                12890: data_o = 32'h00000000 /* 0xc968 */;
                12891: data_o = 32'h00000000 /* 0xc96c */;
                12892: data_o = 32'h00000000 /* 0xc970 */;
                12893: data_o = 32'h00000000 /* 0xc974 */;
                12894: data_o = 32'h00000000 /* 0xc978 */;
                12895: data_o = 32'h00000000 /* 0xc97c */;
                12896: data_o = 32'h00000000 /* 0xc980 */;
                12897: data_o = 32'h00000000 /* 0xc984 */;
                12898: data_o = 32'h00000000 /* 0xc988 */;
                12899: data_o = 32'h00000000 /* 0xc98c */;
                12900: data_o = 32'h00000000 /* 0xc990 */;
                12901: data_o = 32'h00000000 /* 0xc994 */;
                12902: data_o = 32'h00000000 /* 0xc998 */;
                12903: data_o = 32'h00000000 /* 0xc99c */;
                12904: data_o = 32'h00000000 /* 0xc9a0 */;
                12905: data_o = 32'h00000000 /* 0xc9a4 */;
                12906: data_o = 32'h00000000 /* 0xc9a8 */;
                12907: data_o = 32'h00000000 /* 0xc9ac */;
                12908: data_o = 32'h00000000 /* 0xc9b0 */;
                12909: data_o = 32'h00000000 /* 0xc9b4 */;
                12910: data_o = 32'h00000000 /* 0xc9b8 */;
                12911: data_o = 32'h00000000 /* 0xc9bc */;
                12912: data_o = 32'h00000000 /* 0xc9c0 */;
                12913: data_o = 32'h00000000 /* 0xc9c4 */;
                12914: data_o = 32'h00000000 /* 0xc9c8 */;
                12915: data_o = 32'h00000000 /* 0xc9cc */;
                12916: data_o = 32'h00000000 /* 0xc9d0 */;
                12917: data_o = 32'h00000000 /* 0xc9d4 */;
                12918: data_o = 32'h00000000 /* 0xc9d8 */;
                12919: data_o = 32'h00000000 /* 0xc9dc */;
                12920: data_o = 32'h00000000 /* 0xc9e0 */;
                12921: data_o = 32'h00000000 /* 0xc9e4 */;
                12922: data_o = 32'h00000000 /* 0xc9e8 */;
                12923: data_o = 32'h00000000 /* 0xc9ec */;
                12924: data_o = 32'h00000000 /* 0xc9f0 */;
                12925: data_o = 32'h00000000 /* 0xc9f4 */;
                12926: data_o = 32'h00000000 /* 0xc9f8 */;
                12927: data_o = 32'h00000000 /* 0xc9fc */;
                12928: data_o = 32'h00000000 /* 0xca00 */;
                12929: data_o = 32'h00000000 /* 0xca04 */;
                12930: data_o = 32'h00000000 /* 0xca08 */;
                12931: data_o = 32'h00000000 /* 0xca0c */;
                12932: data_o = 32'h00000000 /* 0xca10 */;
                12933: data_o = 32'h00000000 /* 0xca14 */;
                12934: data_o = 32'h00000000 /* 0xca18 */;
                12935: data_o = 32'h00000000 /* 0xca1c */;
                12936: data_o = 32'h00000000 /* 0xca20 */;
                12937: data_o = 32'h00000000 /* 0xca24 */;
                12938: data_o = 32'h00000000 /* 0xca28 */;
                12939: data_o = 32'h00000000 /* 0xca2c */;
                12940: data_o = 32'h00000000 /* 0xca30 */;
                12941: data_o = 32'h00000000 /* 0xca34 */;
                12942: data_o = 32'h00000000 /* 0xca38 */;
                12943: data_o = 32'h00000000 /* 0xca3c */;
                12944: data_o = 32'h00000000 /* 0xca40 */;
                12945: data_o = 32'h00000000 /* 0xca44 */;
                12946: data_o = 32'h00000000 /* 0xca48 */;
                12947: data_o = 32'h00000000 /* 0xca4c */;
                12948: data_o = 32'h00000000 /* 0xca50 */;
                12949: data_o = 32'h00000000 /* 0xca54 */;
                12950: data_o = 32'h00000000 /* 0xca58 */;
                12951: data_o = 32'h00000000 /* 0xca5c */;
                12952: data_o = 32'h00000000 /* 0xca60 */;
                12953: data_o = 32'h00000000 /* 0xca64 */;
                12954: data_o = 32'h00000000 /* 0xca68 */;
                12955: data_o = 32'h00000000 /* 0xca6c */;
                12956: data_o = 32'h00000000 /* 0xca70 */;
                12957: data_o = 32'h00000000 /* 0xca74 */;
                12958: data_o = 32'h00000000 /* 0xca78 */;
                12959: data_o = 32'h00000000 /* 0xca7c */;
                12960: data_o = 32'h00000000 /* 0xca80 */;
                12961: data_o = 32'h00000000 /* 0xca84 */;
                12962: data_o = 32'h00000000 /* 0xca88 */;
                12963: data_o = 32'h00000000 /* 0xca8c */;
                12964: data_o = 32'h00000000 /* 0xca90 */;
                12965: data_o = 32'h00000000 /* 0xca94 */;
                12966: data_o = 32'h00000000 /* 0xca98 */;
                12967: data_o = 32'h00000000 /* 0xca9c */;
                12968: data_o = 32'h00000000 /* 0xcaa0 */;
                12969: data_o = 32'h00000000 /* 0xcaa4 */;
                12970: data_o = 32'h00000000 /* 0xcaa8 */;
                12971: data_o = 32'h00000000 /* 0xcaac */;
                12972: data_o = 32'h00000000 /* 0xcab0 */;
                12973: data_o = 32'h00000000 /* 0xcab4 */;
                12974: data_o = 32'h00000000 /* 0xcab8 */;
                12975: data_o = 32'h00000000 /* 0xcabc */;
                12976: data_o = 32'h00000000 /* 0xcac0 */;
                12977: data_o = 32'h00000000 /* 0xcac4 */;
                12978: data_o = 32'h00000000 /* 0xcac8 */;
                12979: data_o = 32'h00000000 /* 0xcacc */;
                12980: data_o = 32'h00000000 /* 0xcad0 */;
                12981: data_o = 32'h00000000 /* 0xcad4 */;
                12982: data_o = 32'h00000000 /* 0xcad8 */;
                12983: data_o = 32'h00000000 /* 0xcadc */;
                12984: data_o = 32'h00000000 /* 0xcae0 */;
                12985: data_o = 32'h00000000 /* 0xcae4 */;
                12986: data_o = 32'h00000000 /* 0xcae8 */;
                12987: data_o = 32'h00000000 /* 0xcaec */;
                12988: data_o = 32'h00000000 /* 0xcaf0 */;
                12989: data_o = 32'h00000000 /* 0xcaf4 */;
                12990: data_o = 32'h00000000 /* 0xcaf8 */;
                12991: data_o = 32'h00000000 /* 0xcafc */;
                12992: data_o = 32'h00000000 /* 0xcb00 */;
                12993: data_o = 32'h00000000 /* 0xcb04 */;
                12994: data_o = 32'h00000000 /* 0xcb08 */;
                12995: data_o = 32'h00000000 /* 0xcb0c */;
                12996: data_o = 32'h00000000 /* 0xcb10 */;
                12997: data_o = 32'h00000000 /* 0xcb14 */;
                12998: data_o = 32'h00000000 /* 0xcb18 */;
                12999: data_o = 32'h00000000 /* 0xcb1c */;
                13000: data_o = 32'h00000000 /* 0xcb20 */;
                13001: data_o = 32'h00000000 /* 0xcb24 */;
                13002: data_o = 32'h00000000 /* 0xcb28 */;
                13003: data_o = 32'h00000000 /* 0xcb2c */;
                13004: data_o = 32'h00000000 /* 0xcb30 */;
                13005: data_o = 32'h00000000 /* 0xcb34 */;
                13006: data_o = 32'h00000000 /* 0xcb38 */;
                13007: data_o = 32'h00000000 /* 0xcb3c */;
                13008: data_o = 32'h00000000 /* 0xcb40 */;
                13009: data_o = 32'h00000000 /* 0xcb44 */;
                13010: data_o = 32'h00000000 /* 0xcb48 */;
                13011: data_o = 32'h00000000 /* 0xcb4c */;
                13012: data_o = 32'h00000000 /* 0xcb50 */;
                13013: data_o = 32'h00000000 /* 0xcb54 */;
                13014: data_o = 32'h00000000 /* 0xcb58 */;
                13015: data_o = 32'h00000000 /* 0xcb5c */;
                13016: data_o = 32'h00000000 /* 0xcb60 */;
                13017: data_o = 32'h00000000 /* 0xcb64 */;
                13018: data_o = 32'h00000000 /* 0xcb68 */;
                13019: data_o = 32'h00000000 /* 0xcb6c */;
                13020: data_o = 32'h00000000 /* 0xcb70 */;
                13021: data_o = 32'h00000000 /* 0xcb74 */;
                13022: data_o = 32'h00000000 /* 0xcb78 */;
                13023: data_o = 32'h00000000 /* 0xcb7c */;
                13024: data_o = 32'h00000000 /* 0xcb80 */;
                13025: data_o = 32'h00000000 /* 0xcb84 */;
                13026: data_o = 32'h00000000 /* 0xcb88 */;
                13027: data_o = 32'h00000000 /* 0xcb8c */;
                13028: data_o = 32'h00000000 /* 0xcb90 */;
                13029: data_o = 32'h00000000 /* 0xcb94 */;
                13030: data_o = 32'h00000000 /* 0xcb98 */;
                13031: data_o = 32'h00000000 /* 0xcb9c */;
                13032: data_o = 32'h00000000 /* 0xcba0 */;
                13033: data_o = 32'h00000000 /* 0xcba4 */;
                13034: data_o = 32'h00000000 /* 0xcba8 */;
                13035: data_o = 32'h00000000 /* 0xcbac */;
                13036: data_o = 32'h00000000 /* 0xcbb0 */;
                13037: data_o = 32'h00000000 /* 0xcbb4 */;
                13038: data_o = 32'h00000000 /* 0xcbb8 */;
                13039: data_o = 32'h00000000 /* 0xcbbc */;
                13040: data_o = 32'h00000000 /* 0xcbc0 */;
                13041: data_o = 32'h00000000 /* 0xcbc4 */;
                13042: data_o = 32'h00000000 /* 0xcbc8 */;
                13043: data_o = 32'h00000000 /* 0xcbcc */;
                13044: data_o = 32'h00000000 /* 0xcbd0 */;
                13045: data_o = 32'h00000000 /* 0xcbd4 */;
                13046: data_o = 32'h00000000 /* 0xcbd8 */;
                13047: data_o = 32'h00000000 /* 0xcbdc */;
                13048: data_o = 32'h00000000 /* 0xcbe0 */;
                13049: data_o = 32'h00000000 /* 0xcbe4 */;
                13050: data_o = 32'h00000000 /* 0xcbe8 */;
                13051: data_o = 32'h00000000 /* 0xcbec */;
                13052: data_o = 32'h00000000 /* 0xcbf0 */;
                13053: data_o = 32'h00000000 /* 0xcbf4 */;
                13054: data_o = 32'h00000000 /* 0xcbf8 */;
                13055: data_o = 32'h00000000 /* 0xcbfc */;
                13056: data_o = 32'h00000000 /* 0xcc00 */;
                13057: data_o = 32'h00000000 /* 0xcc04 */;
                13058: data_o = 32'h00000000 /* 0xcc08 */;
                13059: data_o = 32'h00000000 /* 0xcc0c */;
                13060: data_o = 32'h00000000 /* 0xcc10 */;
                13061: data_o = 32'h00000000 /* 0xcc14 */;
                13062: data_o = 32'h00000000 /* 0xcc18 */;
                13063: data_o = 32'h00000000 /* 0xcc1c */;
                13064: data_o = 32'h00000000 /* 0xcc20 */;
                13065: data_o = 32'h00000000 /* 0xcc24 */;
                13066: data_o = 32'h00000000 /* 0xcc28 */;
                13067: data_o = 32'h00000000 /* 0xcc2c */;
                13068: data_o = 32'h00000000 /* 0xcc30 */;
                13069: data_o = 32'h00000000 /* 0xcc34 */;
                13070: data_o = 32'h00000000 /* 0xcc38 */;
                13071: data_o = 32'h00000000 /* 0xcc3c */;
                13072: data_o = 32'h00000000 /* 0xcc40 */;
                13073: data_o = 32'h00000000 /* 0xcc44 */;
                13074: data_o = 32'h00000000 /* 0xcc48 */;
                13075: data_o = 32'h00000000 /* 0xcc4c */;
                13076: data_o = 32'h00000000 /* 0xcc50 */;
                13077: data_o = 32'h00000000 /* 0xcc54 */;
                13078: data_o = 32'h00000000 /* 0xcc58 */;
                13079: data_o = 32'h00000000 /* 0xcc5c */;
                13080: data_o = 32'h00000000 /* 0xcc60 */;
                13081: data_o = 32'h00000000 /* 0xcc64 */;
                13082: data_o = 32'h00000000 /* 0xcc68 */;
                13083: data_o = 32'h00000000 /* 0xcc6c */;
                13084: data_o = 32'h00000000 /* 0xcc70 */;
                13085: data_o = 32'h00000000 /* 0xcc74 */;
                13086: data_o = 32'h00000000 /* 0xcc78 */;
                13087: data_o = 32'h00000000 /* 0xcc7c */;
                13088: data_o = 32'h00000000 /* 0xcc80 */;
                13089: data_o = 32'h00000000 /* 0xcc84 */;
                13090: data_o = 32'h00000000 /* 0xcc88 */;
                13091: data_o = 32'h00000000 /* 0xcc8c */;
                13092: data_o = 32'h00000000 /* 0xcc90 */;
                13093: data_o = 32'h00000000 /* 0xcc94 */;
                13094: data_o = 32'h00000000 /* 0xcc98 */;
                13095: data_o = 32'h00000000 /* 0xcc9c */;
                13096: data_o = 32'h00000000 /* 0xcca0 */;
                13097: data_o = 32'h00000000 /* 0xcca4 */;
                13098: data_o = 32'h00000000 /* 0xcca8 */;
                13099: data_o = 32'h00000000 /* 0xccac */;
                13100: data_o = 32'h00000000 /* 0xccb0 */;
                13101: data_o = 32'h00000000 /* 0xccb4 */;
                13102: data_o = 32'h00000000 /* 0xccb8 */;
                13103: data_o = 32'h00000000 /* 0xccbc */;
                13104: data_o = 32'h00000000 /* 0xccc0 */;
                13105: data_o = 32'h00000000 /* 0xccc4 */;
                13106: data_o = 32'h00000000 /* 0xccc8 */;
                13107: data_o = 32'h00000000 /* 0xcccc */;
                13108: data_o = 32'h00000000 /* 0xccd0 */;
                13109: data_o = 32'h00000000 /* 0xccd4 */;
                13110: data_o = 32'h00000000 /* 0xccd8 */;
                13111: data_o = 32'h00000000 /* 0xccdc */;
                13112: data_o = 32'h00000000 /* 0xcce0 */;
                13113: data_o = 32'h00000000 /* 0xcce4 */;
                13114: data_o = 32'h00000000 /* 0xcce8 */;
                13115: data_o = 32'h00000000 /* 0xccec */;
                13116: data_o = 32'h00000000 /* 0xccf0 */;
                13117: data_o = 32'h00000000 /* 0xccf4 */;
                13118: data_o = 32'h00000000 /* 0xccf8 */;
                13119: data_o = 32'h00000000 /* 0xccfc */;
                13120: data_o = 32'h00000000 /* 0xcd00 */;
                13121: data_o = 32'h00000000 /* 0xcd04 */;
                13122: data_o = 32'h00000000 /* 0xcd08 */;
                13123: data_o = 32'h00000000 /* 0xcd0c */;
                13124: data_o = 32'h00000000 /* 0xcd10 */;
                13125: data_o = 32'h00000000 /* 0xcd14 */;
                13126: data_o = 32'h00000000 /* 0xcd18 */;
                13127: data_o = 32'h00000000 /* 0xcd1c */;
                13128: data_o = 32'h00000000 /* 0xcd20 */;
                13129: data_o = 32'h00000000 /* 0xcd24 */;
                13130: data_o = 32'h00000000 /* 0xcd28 */;
                13131: data_o = 32'h00000000 /* 0xcd2c */;
                13132: data_o = 32'h00000000 /* 0xcd30 */;
                13133: data_o = 32'h00000000 /* 0xcd34 */;
                13134: data_o = 32'h00000000 /* 0xcd38 */;
                13135: data_o = 32'h00000000 /* 0xcd3c */;
                13136: data_o = 32'h00000000 /* 0xcd40 */;
                13137: data_o = 32'h00000000 /* 0xcd44 */;
                13138: data_o = 32'h00000000 /* 0xcd48 */;
                13139: data_o = 32'h00000000 /* 0xcd4c */;
                13140: data_o = 32'h00000000 /* 0xcd50 */;
                13141: data_o = 32'h00000000 /* 0xcd54 */;
                13142: data_o = 32'h00000000 /* 0xcd58 */;
                13143: data_o = 32'h00000000 /* 0xcd5c */;
                13144: data_o = 32'h00000000 /* 0xcd60 */;
                13145: data_o = 32'h00000000 /* 0xcd64 */;
                13146: data_o = 32'h00000000 /* 0xcd68 */;
                13147: data_o = 32'h00000000 /* 0xcd6c */;
                13148: data_o = 32'h00000000 /* 0xcd70 */;
                13149: data_o = 32'h00000000 /* 0xcd74 */;
                13150: data_o = 32'h00000000 /* 0xcd78 */;
                13151: data_o = 32'h00000000 /* 0xcd7c */;
                13152: data_o = 32'h00000000 /* 0xcd80 */;
                13153: data_o = 32'h00000000 /* 0xcd84 */;
                13154: data_o = 32'h00000000 /* 0xcd88 */;
                13155: data_o = 32'h00000000 /* 0xcd8c */;
                13156: data_o = 32'h00000000 /* 0xcd90 */;
                13157: data_o = 32'h00000000 /* 0xcd94 */;
                13158: data_o = 32'h00000000 /* 0xcd98 */;
                13159: data_o = 32'h00000000 /* 0xcd9c */;
                13160: data_o = 32'h00000000 /* 0xcda0 */;
                13161: data_o = 32'h00000000 /* 0xcda4 */;
                13162: data_o = 32'h00000000 /* 0xcda8 */;
                13163: data_o = 32'h00000000 /* 0xcdac */;
                13164: data_o = 32'h00000000 /* 0xcdb0 */;
                13165: data_o = 32'h00000000 /* 0xcdb4 */;
                13166: data_o = 32'h00000000 /* 0xcdb8 */;
                13167: data_o = 32'h00000000 /* 0xcdbc */;
                13168: data_o = 32'h00000000 /* 0xcdc0 */;
                13169: data_o = 32'h00000000 /* 0xcdc4 */;
                13170: data_o = 32'h00000000 /* 0xcdc8 */;
                13171: data_o = 32'h00000000 /* 0xcdcc */;
                13172: data_o = 32'h00000000 /* 0xcdd0 */;
                13173: data_o = 32'h00000000 /* 0xcdd4 */;
                13174: data_o = 32'h00000000 /* 0xcdd8 */;
                13175: data_o = 32'h00000000 /* 0xcddc */;
                13176: data_o = 32'h00000000 /* 0xcde0 */;
                13177: data_o = 32'h00000000 /* 0xcde4 */;
                13178: data_o = 32'h00000000 /* 0xcde8 */;
                13179: data_o = 32'h00000000 /* 0xcdec */;
                13180: data_o = 32'h00000000 /* 0xcdf0 */;
                13181: data_o = 32'h00000000 /* 0xcdf4 */;
                13182: data_o = 32'h00000000 /* 0xcdf8 */;
                13183: data_o = 32'h00000000 /* 0xcdfc */;
                13184: data_o = 32'h00000000 /* 0xce00 */;
                13185: data_o = 32'h00000000 /* 0xce04 */;
                13186: data_o = 32'h00000000 /* 0xce08 */;
                13187: data_o = 32'h00000000 /* 0xce0c */;
                13188: data_o = 32'h00000000 /* 0xce10 */;
                13189: data_o = 32'h00000000 /* 0xce14 */;
                13190: data_o = 32'h00000000 /* 0xce18 */;
                13191: data_o = 32'h00000000 /* 0xce1c */;
                13192: data_o = 32'h00000000 /* 0xce20 */;
                13193: data_o = 32'h00000000 /* 0xce24 */;
                13194: data_o = 32'h00000000 /* 0xce28 */;
                13195: data_o = 32'h00000000 /* 0xce2c */;
                13196: data_o = 32'h00000000 /* 0xce30 */;
                13197: data_o = 32'h00000000 /* 0xce34 */;
                13198: data_o = 32'h00000000 /* 0xce38 */;
                13199: data_o = 32'h00000000 /* 0xce3c */;
                13200: data_o = 32'h00000000 /* 0xce40 */;
                13201: data_o = 32'h00000000 /* 0xce44 */;
                13202: data_o = 32'h00000000 /* 0xce48 */;
                13203: data_o = 32'h00000000 /* 0xce4c */;
                13204: data_o = 32'h00000000 /* 0xce50 */;
                13205: data_o = 32'h00000000 /* 0xce54 */;
                13206: data_o = 32'h00000000 /* 0xce58 */;
                13207: data_o = 32'h00000000 /* 0xce5c */;
                13208: data_o = 32'h00000000 /* 0xce60 */;
                13209: data_o = 32'h00000000 /* 0xce64 */;
                13210: data_o = 32'h00000000 /* 0xce68 */;
                13211: data_o = 32'h00000000 /* 0xce6c */;
                13212: data_o = 32'h00000000 /* 0xce70 */;
                13213: data_o = 32'h00000000 /* 0xce74 */;
                13214: data_o = 32'h00000000 /* 0xce78 */;
                13215: data_o = 32'h00000000 /* 0xce7c */;
                13216: data_o = 32'h00000000 /* 0xce80 */;
                13217: data_o = 32'h00000000 /* 0xce84 */;
                13218: data_o = 32'h00000000 /* 0xce88 */;
                13219: data_o = 32'h00000000 /* 0xce8c */;
                13220: data_o = 32'h00000000 /* 0xce90 */;
                13221: data_o = 32'h00000000 /* 0xce94 */;
                13222: data_o = 32'h00000000 /* 0xce98 */;
                13223: data_o = 32'h00000000 /* 0xce9c */;
                13224: data_o = 32'h00000000 /* 0xcea0 */;
                13225: data_o = 32'h00000000 /* 0xcea4 */;
                13226: data_o = 32'h00000000 /* 0xcea8 */;
                13227: data_o = 32'h00000000 /* 0xceac */;
                13228: data_o = 32'h00000000 /* 0xceb0 */;
                13229: data_o = 32'h00000000 /* 0xceb4 */;
                13230: data_o = 32'h00000000 /* 0xceb8 */;
                13231: data_o = 32'h00000000 /* 0xcebc */;
                13232: data_o = 32'h00000000 /* 0xcec0 */;
                13233: data_o = 32'h00000000 /* 0xcec4 */;
                13234: data_o = 32'h00000000 /* 0xcec8 */;
                13235: data_o = 32'h00000000 /* 0xcecc */;
                13236: data_o = 32'h00000000 /* 0xced0 */;
                13237: data_o = 32'h00000000 /* 0xced4 */;
                13238: data_o = 32'h00000000 /* 0xced8 */;
                13239: data_o = 32'h00000000 /* 0xcedc */;
                13240: data_o = 32'h00000000 /* 0xcee0 */;
                13241: data_o = 32'h00000000 /* 0xcee4 */;
                13242: data_o = 32'h00000000 /* 0xcee8 */;
                13243: data_o = 32'h00000000 /* 0xceec */;
                13244: data_o = 32'h00000000 /* 0xcef0 */;
                13245: data_o = 32'h00000000 /* 0xcef4 */;
                13246: data_o = 32'h00000000 /* 0xcef8 */;
                13247: data_o = 32'h00000000 /* 0xcefc */;
                13248: data_o = 32'h00000000 /* 0xcf00 */;
                13249: data_o = 32'h00000000 /* 0xcf04 */;
                13250: data_o = 32'h00000000 /* 0xcf08 */;
                13251: data_o = 32'h00000000 /* 0xcf0c */;
                13252: data_o = 32'h00000000 /* 0xcf10 */;
                13253: data_o = 32'h00000000 /* 0xcf14 */;
                13254: data_o = 32'h00000000 /* 0xcf18 */;
                13255: data_o = 32'h00000000 /* 0xcf1c */;
                13256: data_o = 32'h00000000 /* 0xcf20 */;
                13257: data_o = 32'h00000000 /* 0xcf24 */;
                13258: data_o = 32'h00000000 /* 0xcf28 */;
                13259: data_o = 32'h00000000 /* 0xcf2c */;
                13260: data_o = 32'h00000000 /* 0xcf30 */;
                13261: data_o = 32'h00000000 /* 0xcf34 */;
                13262: data_o = 32'h00000000 /* 0xcf38 */;
                13263: data_o = 32'h00000000 /* 0xcf3c */;
                13264: data_o = 32'h00000000 /* 0xcf40 */;
                13265: data_o = 32'h00000000 /* 0xcf44 */;
                13266: data_o = 32'h00000000 /* 0xcf48 */;
                13267: data_o = 32'h00000000 /* 0xcf4c */;
                13268: data_o = 32'h00000000 /* 0xcf50 */;
                13269: data_o = 32'h00000000 /* 0xcf54 */;
                13270: data_o = 32'h00000000 /* 0xcf58 */;
                13271: data_o = 32'h00000000 /* 0xcf5c */;
                13272: data_o = 32'h00000000 /* 0xcf60 */;
                13273: data_o = 32'h00000000 /* 0xcf64 */;
                13274: data_o = 32'h00000000 /* 0xcf68 */;
                13275: data_o = 32'h00000000 /* 0xcf6c */;
                13276: data_o = 32'h00000000 /* 0xcf70 */;
                13277: data_o = 32'h00000000 /* 0xcf74 */;
                13278: data_o = 32'h00000000 /* 0xcf78 */;
                13279: data_o = 32'h00000000 /* 0xcf7c */;
                13280: data_o = 32'h00000000 /* 0xcf80 */;
                13281: data_o = 32'h00000000 /* 0xcf84 */;
                13282: data_o = 32'h00000000 /* 0xcf88 */;
                13283: data_o = 32'h00000000 /* 0xcf8c */;
                13284: data_o = 32'h00000000 /* 0xcf90 */;
                13285: data_o = 32'h00000000 /* 0xcf94 */;
                13286: data_o = 32'h00000000 /* 0xcf98 */;
                13287: data_o = 32'h00000000 /* 0xcf9c */;
                13288: data_o = 32'h00000000 /* 0xcfa0 */;
                13289: data_o = 32'h00000000 /* 0xcfa4 */;
                13290: data_o = 32'h00000000 /* 0xcfa8 */;
                13291: data_o = 32'h00000000 /* 0xcfac */;
                13292: data_o = 32'h00000000 /* 0xcfb0 */;
                13293: data_o = 32'h00000000 /* 0xcfb4 */;
                13294: data_o = 32'h00000000 /* 0xcfb8 */;
                13295: data_o = 32'h00000000 /* 0xcfbc */;
                13296: data_o = 32'h00000000 /* 0xcfc0 */;
                13297: data_o = 32'h00000000 /* 0xcfc4 */;
                13298: data_o = 32'h00000000 /* 0xcfc8 */;
                13299: data_o = 32'h00000000 /* 0xcfcc */;
                13300: data_o = 32'h00000000 /* 0xcfd0 */;
                13301: data_o = 32'h00000000 /* 0xcfd4 */;
                13302: data_o = 32'h00000000 /* 0xcfd8 */;
                13303: data_o = 32'h00000000 /* 0xcfdc */;
                13304: data_o = 32'h00000000 /* 0xcfe0 */;
                13305: data_o = 32'h00000000 /* 0xcfe4 */;
                13306: data_o = 32'h00000000 /* 0xcfe8 */;
                13307: data_o = 32'h00000000 /* 0xcfec */;
                13308: data_o = 32'h00000000 /* 0xcff0 */;
                13309: data_o = 32'h00000000 /* 0xcff4 */;
                13310: data_o = 32'h00000000 /* 0xcff8 */;
                13311: data_o = 32'h00000000 /* 0xcffc */;
                13312: data_o = 32'h00000000 /* 0xd000 */;
                13313: data_o = 32'h00000000 /* 0xd004 */;
                13314: data_o = 32'h00000000 /* 0xd008 */;
                13315: data_o = 32'h00000000 /* 0xd00c */;
                13316: data_o = 32'h00000000 /* 0xd010 */;
                13317: data_o = 32'h00000000 /* 0xd014 */;
                13318: data_o = 32'h00000000 /* 0xd018 */;
                13319: data_o = 32'h00000000 /* 0xd01c */;
                13320: data_o = 32'h00000000 /* 0xd020 */;
                13321: data_o = 32'h00000000 /* 0xd024 */;
                13322: data_o = 32'h00000000 /* 0xd028 */;
                13323: data_o = 32'h00000000 /* 0xd02c */;
                13324: data_o = 32'h00000000 /* 0xd030 */;
                13325: data_o = 32'h00000000 /* 0xd034 */;
                13326: data_o = 32'h00000000 /* 0xd038 */;
                13327: data_o = 32'h00000000 /* 0xd03c */;
                13328: data_o = 32'h00000000 /* 0xd040 */;
                13329: data_o = 32'h00000000 /* 0xd044 */;
                13330: data_o = 32'h00000000 /* 0xd048 */;
                13331: data_o = 32'h00000000 /* 0xd04c */;
                13332: data_o = 32'h00000000 /* 0xd050 */;
                13333: data_o = 32'h00000000 /* 0xd054 */;
                13334: data_o = 32'h00000000 /* 0xd058 */;
                13335: data_o = 32'h00000000 /* 0xd05c */;
                13336: data_o = 32'h00000000 /* 0xd060 */;
                13337: data_o = 32'h00000000 /* 0xd064 */;
                13338: data_o = 32'h00000000 /* 0xd068 */;
                13339: data_o = 32'h00000000 /* 0xd06c */;
                13340: data_o = 32'h00000000 /* 0xd070 */;
                13341: data_o = 32'h00000000 /* 0xd074 */;
                13342: data_o = 32'h00000000 /* 0xd078 */;
                13343: data_o = 32'h00000000 /* 0xd07c */;
                13344: data_o = 32'h00000000 /* 0xd080 */;
                13345: data_o = 32'h00000000 /* 0xd084 */;
                13346: data_o = 32'h00000000 /* 0xd088 */;
                13347: data_o = 32'h00000000 /* 0xd08c */;
                13348: data_o = 32'h00000000 /* 0xd090 */;
                13349: data_o = 32'h00000000 /* 0xd094 */;
                13350: data_o = 32'h00000000 /* 0xd098 */;
                13351: data_o = 32'h00000000 /* 0xd09c */;
                13352: data_o = 32'h00000000 /* 0xd0a0 */;
                13353: data_o = 32'h00000000 /* 0xd0a4 */;
                13354: data_o = 32'h00000000 /* 0xd0a8 */;
                13355: data_o = 32'h00000000 /* 0xd0ac */;
                13356: data_o = 32'h00000000 /* 0xd0b0 */;
                13357: data_o = 32'h00000000 /* 0xd0b4 */;
                13358: data_o = 32'h00000000 /* 0xd0b8 */;
                13359: data_o = 32'h00000000 /* 0xd0bc */;
                13360: data_o = 32'h00000000 /* 0xd0c0 */;
                13361: data_o = 32'h00000000 /* 0xd0c4 */;
                13362: data_o = 32'h00000000 /* 0xd0c8 */;
                13363: data_o = 32'h00000000 /* 0xd0cc */;
                13364: data_o = 32'h00000000 /* 0xd0d0 */;
                13365: data_o = 32'h00000000 /* 0xd0d4 */;
                13366: data_o = 32'h00000000 /* 0xd0d8 */;
                13367: data_o = 32'h00000000 /* 0xd0dc */;
                13368: data_o = 32'h00000000 /* 0xd0e0 */;
                13369: data_o = 32'h00000000 /* 0xd0e4 */;
                13370: data_o = 32'h00000000 /* 0xd0e8 */;
                13371: data_o = 32'h00000000 /* 0xd0ec */;
                13372: data_o = 32'h00000000 /* 0xd0f0 */;
                13373: data_o = 32'h00000000 /* 0xd0f4 */;
                13374: data_o = 32'h00000000 /* 0xd0f8 */;
                13375: data_o = 32'h00000000 /* 0xd0fc */;
                13376: data_o = 32'h00000000 /* 0xd100 */;
                13377: data_o = 32'h00000000 /* 0xd104 */;
                13378: data_o = 32'h00000000 /* 0xd108 */;
                13379: data_o = 32'h00000000 /* 0xd10c */;
                13380: data_o = 32'h00000000 /* 0xd110 */;
                13381: data_o = 32'h00000000 /* 0xd114 */;
                13382: data_o = 32'h00000000 /* 0xd118 */;
                13383: data_o = 32'h00000000 /* 0xd11c */;
                13384: data_o = 32'h00000000 /* 0xd120 */;
                13385: data_o = 32'h00000000 /* 0xd124 */;
                13386: data_o = 32'h00000000 /* 0xd128 */;
                13387: data_o = 32'h00000000 /* 0xd12c */;
                13388: data_o = 32'h00000000 /* 0xd130 */;
                13389: data_o = 32'h00000000 /* 0xd134 */;
                13390: data_o = 32'h00000000 /* 0xd138 */;
                13391: data_o = 32'h00000000 /* 0xd13c */;
                13392: data_o = 32'h00000000 /* 0xd140 */;
                13393: data_o = 32'h00000000 /* 0xd144 */;
                13394: data_o = 32'h00000000 /* 0xd148 */;
                13395: data_o = 32'h00000000 /* 0xd14c */;
                13396: data_o = 32'h00000000 /* 0xd150 */;
                13397: data_o = 32'h00000000 /* 0xd154 */;
                13398: data_o = 32'h00000000 /* 0xd158 */;
                13399: data_o = 32'h00000000 /* 0xd15c */;
                13400: data_o = 32'h00000000 /* 0xd160 */;
                13401: data_o = 32'h00000000 /* 0xd164 */;
                13402: data_o = 32'h00000000 /* 0xd168 */;
                13403: data_o = 32'h00000000 /* 0xd16c */;
                13404: data_o = 32'h00000000 /* 0xd170 */;
                13405: data_o = 32'h00000000 /* 0xd174 */;
                13406: data_o = 32'h00000000 /* 0xd178 */;
                13407: data_o = 32'h00000000 /* 0xd17c */;
                13408: data_o = 32'h00000000 /* 0xd180 */;
                13409: data_o = 32'h00000000 /* 0xd184 */;
                13410: data_o = 32'h00000000 /* 0xd188 */;
                13411: data_o = 32'h00000000 /* 0xd18c */;
                13412: data_o = 32'h00000000 /* 0xd190 */;
                13413: data_o = 32'h00000000 /* 0xd194 */;
                13414: data_o = 32'h00000000 /* 0xd198 */;
                13415: data_o = 32'h00000000 /* 0xd19c */;
                13416: data_o = 32'h00000000 /* 0xd1a0 */;
                13417: data_o = 32'h00000000 /* 0xd1a4 */;
                13418: data_o = 32'h00000000 /* 0xd1a8 */;
                13419: data_o = 32'h00000000 /* 0xd1ac */;
                13420: data_o = 32'h00000000 /* 0xd1b0 */;
                13421: data_o = 32'h00000000 /* 0xd1b4 */;
                13422: data_o = 32'h00000000 /* 0xd1b8 */;
                13423: data_o = 32'h00000000 /* 0xd1bc */;
                13424: data_o = 32'h00000000 /* 0xd1c0 */;
                13425: data_o = 32'h00000000 /* 0xd1c4 */;
                13426: data_o = 32'h00000000 /* 0xd1c8 */;
                13427: data_o = 32'h00000000 /* 0xd1cc */;
                13428: data_o = 32'h00000000 /* 0xd1d0 */;
                13429: data_o = 32'h00000000 /* 0xd1d4 */;
                13430: data_o = 32'h00000000 /* 0xd1d8 */;
                13431: data_o = 32'h00000000 /* 0xd1dc */;
                13432: data_o = 32'h00000000 /* 0xd1e0 */;
                13433: data_o = 32'h00000000 /* 0xd1e4 */;
                13434: data_o = 32'h00000000 /* 0xd1e8 */;
                13435: data_o = 32'h00000000 /* 0xd1ec */;
                13436: data_o = 32'h00000000 /* 0xd1f0 */;
                13437: data_o = 32'h00000000 /* 0xd1f4 */;
                13438: data_o = 32'h00000000 /* 0xd1f8 */;
                13439: data_o = 32'h00000000 /* 0xd1fc */;
                13440: data_o = 32'h00000000 /* 0xd200 */;
                13441: data_o = 32'h00000000 /* 0xd204 */;
                13442: data_o = 32'h00000000 /* 0xd208 */;
                13443: data_o = 32'h00000000 /* 0xd20c */;
                13444: data_o = 32'h00000000 /* 0xd210 */;
                13445: data_o = 32'h00000000 /* 0xd214 */;
                13446: data_o = 32'h00000000 /* 0xd218 */;
                13447: data_o = 32'h00000000 /* 0xd21c */;
                13448: data_o = 32'h00000000 /* 0xd220 */;
                13449: data_o = 32'h00000000 /* 0xd224 */;
                13450: data_o = 32'h00000000 /* 0xd228 */;
                13451: data_o = 32'h00000000 /* 0xd22c */;
                13452: data_o = 32'h00000000 /* 0xd230 */;
                13453: data_o = 32'h00000000 /* 0xd234 */;
                13454: data_o = 32'h00000000 /* 0xd238 */;
                13455: data_o = 32'h00000000 /* 0xd23c */;
                13456: data_o = 32'h00000000 /* 0xd240 */;
                13457: data_o = 32'h00000000 /* 0xd244 */;
                13458: data_o = 32'h00000000 /* 0xd248 */;
                13459: data_o = 32'h00000000 /* 0xd24c */;
                13460: data_o = 32'h00000000 /* 0xd250 */;
                13461: data_o = 32'h00000000 /* 0xd254 */;
                13462: data_o = 32'h00000000 /* 0xd258 */;
                13463: data_o = 32'h00000000 /* 0xd25c */;
                13464: data_o = 32'h00000000 /* 0xd260 */;
                13465: data_o = 32'h00000000 /* 0xd264 */;
                13466: data_o = 32'h00000000 /* 0xd268 */;
                13467: data_o = 32'h00000000 /* 0xd26c */;
                13468: data_o = 32'h00000000 /* 0xd270 */;
                13469: data_o = 32'h00000000 /* 0xd274 */;
                13470: data_o = 32'h00000000 /* 0xd278 */;
                13471: data_o = 32'h00000000 /* 0xd27c */;
                13472: data_o = 32'h00000000 /* 0xd280 */;
                13473: data_o = 32'h00000000 /* 0xd284 */;
                13474: data_o = 32'h00000000 /* 0xd288 */;
                13475: data_o = 32'h00000000 /* 0xd28c */;
                13476: data_o = 32'h00000000 /* 0xd290 */;
                13477: data_o = 32'h00000000 /* 0xd294 */;
                13478: data_o = 32'h00000000 /* 0xd298 */;
                13479: data_o = 32'h00000000 /* 0xd29c */;
                13480: data_o = 32'h00000000 /* 0xd2a0 */;
                13481: data_o = 32'h00000000 /* 0xd2a4 */;
                13482: data_o = 32'h00000000 /* 0xd2a8 */;
                13483: data_o = 32'h00000000 /* 0xd2ac */;
                13484: data_o = 32'h00000000 /* 0xd2b0 */;
                13485: data_o = 32'h00000000 /* 0xd2b4 */;
                13486: data_o = 32'h00000000 /* 0xd2b8 */;
                13487: data_o = 32'h00000000 /* 0xd2bc */;
                13488: data_o = 32'h00000000 /* 0xd2c0 */;
                13489: data_o = 32'h00000000 /* 0xd2c4 */;
                13490: data_o = 32'h00000000 /* 0xd2c8 */;
                13491: data_o = 32'h00000000 /* 0xd2cc */;
                13492: data_o = 32'h00000000 /* 0xd2d0 */;
                13493: data_o = 32'h00000000 /* 0xd2d4 */;
                13494: data_o = 32'h00000000 /* 0xd2d8 */;
                13495: data_o = 32'h00000000 /* 0xd2dc */;
                13496: data_o = 32'h00000000 /* 0xd2e0 */;
                13497: data_o = 32'h00000000 /* 0xd2e4 */;
                13498: data_o = 32'h00000000 /* 0xd2e8 */;
                13499: data_o = 32'h00000000 /* 0xd2ec */;
                13500: data_o = 32'h00000000 /* 0xd2f0 */;
                13501: data_o = 32'h00000000 /* 0xd2f4 */;
                13502: data_o = 32'h00000000 /* 0xd2f8 */;
                13503: data_o = 32'h00000000 /* 0xd2fc */;
                13504: data_o = 32'h00000000 /* 0xd300 */;
                13505: data_o = 32'h00000000 /* 0xd304 */;
                13506: data_o = 32'h00000000 /* 0xd308 */;
                13507: data_o = 32'h00000000 /* 0xd30c */;
                13508: data_o = 32'h00000000 /* 0xd310 */;
                13509: data_o = 32'h00000000 /* 0xd314 */;
                13510: data_o = 32'h00000000 /* 0xd318 */;
                13511: data_o = 32'h00000000 /* 0xd31c */;
                13512: data_o = 32'h00000000 /* 0xd320 */;
                13513: data_o = 32'h00000000 /* 0xd324 */;
                13514: data_o = 32'h00000000 /* 0xd328 */;
                13515: data_o = 32'h00000000 /* 0xd32c */;
                13516: data_o = 32'h00000000 /* 0xd330 */;
                13517: data_o = 32'h00000000 /* 0xd334 */;
                13518: data_o = 32'h00000000 /* 0xd338 */;
                13519: data_o = 32'h00000000 /* 0xd33c */;
                13520: data_o = 32'h00000000 /* 0xd340 */;
                13521: data_o = 32'h00000000 /* 0xd344 */;
                13522: data_o = 32'h00000000 /* 0xd348 */;
                13523: data_o = 32'h00000000 /* 0xd34c */;
                13524: data_o = 32'h00000000 /* 0xd350 */;
                13525: data_o = 32'h00000000 /* 0xd354 */;
                13526: data_o = 32'h00000000 /* 0xd358 */;
                13527: data_o = 32'h00000000 /* 0xd35c */;
                13528: data_o = 32'h00000000 /* 0xd360 */;
                13529: data_o = 32'h00000000 /* 0xd364 */;
                13530: data_o = 32'h00000000 /* 0xd368 */;
                13531: data_o = 32'h00000000 /* 0xd36c */;
                13532: data_o = 32'h00000000 /* 0xd370 */;
                13533: data_o = 32'h00000000 /* 0xd374 */;
                13534: data_o = 32'h00000000 /* 0xd378 */;
                13535: data_o = 32'h00000000 /* 0xd37c */;
                13536: data_o = 32'h00000000 /* 0xd380 */;
                13537: data_o = 32'h00000000 /* 0xd384 */;
                13538: data_o = 32'h00000000 /* 0xd388 */;
                13539: data_o = 32'h00000000 /* 0xd38c */;
                13540: data_o = 32'h00000000 /* 0xd390 */;
                13541: data_o = 32'h00000000 /* 0xd394 */;
                13542: data_o = 32'h00000000 /* 0xd398 */;
                13543: data_o = 32'h00000000 /* 0xd39c */;
                13544: data_o = 32'h00000000 /* 0xd3a0 */;
                13545: data_o = 32'h00000000 /* 0xd3a4 */;
                13546: data_o = 32'h00000000 /* 0xd3a8 */;
                13547: data_o = 32'h00000000 /* 0xd3ac */;
                13548: data_o = 32'h00000000 /* 0xd3b0 */;
                13549: data_o = 32'h00000000 /* 0xd3b4 */;
                13550: data_o = 32'h00000000 /* 0xd3b8 */;
                13551: data_o = 32'h00000000 /* 0xd3bc */;
                13552: data_o = 32'h00000000 /* 0xd3c0 */;
                13553: data_o = 32'h00000000 /* 0xd3c4 */;
                13554: data_o = 32'h00000000 /* 0xd3c8 */;
                13555: data_o = 32'h00000000 /* 0xd3cc */;
                13556: data_o = 32'h00000000 /* 0xd3d0 */;
                13557: data_o = 32'h00000000 /* 0xd3d4 */;
                13558: data_o = 32'h00000000 /* 0xd3d8 */;
                13559: data_o = 32'h00000000 /* 0xd3dc */;
                13560: data_o = 32'h00000000 /* 0xd3e0 */;
                13561: data_o = 32'h00000000 /* 0xd3e4 */;
                13562: data_o = 32'h00000000 /* 0xd3e8 */;
                13563: data_o = 32'h00000000 /* 0xd3ec */;
                13564: data_o = 32'h00000000 /* 0xd3f0 */;
                13565: data_o = 32'h00000000 /* 0xd3f4 */;
                13566: data_o = 32'h00000000 /* 0xd3f8 */;
                13567: data_o = 32'h00000000 /* 0xd3fc */;
                13568: data_o = 32'h00000000 /* 0xd400 */;
                13569: data_o = 32'h00000000 /* 0xd404 */;
                13570: data_o = 32'h00000000 /* 0xd408 */;
                13571: data_o = 32'h00000000 /* 0xd40c */;
                13572: data_o = 32'h00000000 /* 0xd410 */;
                13573: data_o = 32'h00000000 /* 0xd414 */;
                13574: data_o = 32'h00000000 /* 0xd418 */;
                13575: data_o = 32'h00000000 /* 0xd41c */;
                13576: data_o = 32'h00000000 /* 0xd420 */;
                13577: data_o = 32'h00000000 /* 0xd424 */;
                13578: data_o = 32'h00000000 /* 0xd428 */;
                13579: data_o = 32'h00000000 /* 0xd42c */;
                13580: data_o = 32'h00000000 /* 0xd430 */;
                13581: data_o = 32'h00000000 /* 0xd434 */;
                13582: data_o = 32'h00000000 /* 0xd438 */;
                13583: data_o = 32'h00000000 /* 0xd43c */;
                13584: data_o = 32'h00000000 /* 0xd440 */;
                13585: data_o = 32'h00000000 /* 0xd444 */;
                13586: data_o = 32'h00000000 /* 0xd448 */;
                13587: data_o = 32'h00000000 /* 0xd44c */;
                13588: data_o = 32'h00000000 /* 0xd450 */;
                13589: data_o = 32'h00000000 /* 0xd454 */;
                13590: data_o = 32'h00000000 /* 0xd458 */;
                13591: data_o = 32'h00000000 /* 0xd45c */;
                13592: data_o = 32'h00000000 /* 0xd460 */;
                13593: data_o = 32'h00000000 /* 0xd464 */;
                13594: data_o = 32'h00000000 /* 0xd468 */;
                13595: data_o = 32'h00000000 /* 0xd46c */;
                13596: data_o = 32'h00000000 /* 0xd470 */;
                13597: data_o = 32'h00000000 /* 0xd474 */;
                13598: data_o = 32'h00000000 /* 0xd478 */;
                13599: data_o = 32'h00000000 /* 0xd47c */;
                13600: data_o = 32'h00000000 /* 0xd480 */;
                13601: data_o = 32'h00000000 /* 0xd484 */;
                13602: data_o = 32'h00000000 /* 0xd488 */;
                13603: data_o = 32'h00000000 /* 0xd48c */;
                13604: data_o = 32'h00000000 /* 0xd490 */;
                13605: data_o = 32'h00000000 /* 0xd494 */;
                13606: data_o = 32'h00000000 /* 0xd498 */;
                13607: data_o = 32'h00000000 /* 0xd49c */;
                13608: data_o = 32'h00000000 /* 0xd4a0 */;
                13609: data_o = 32'h00000000 /* 0xd4a4 */;
                13610: data_o = 32'h00000000 /* 0xd4a8 */;
                13611: data_o = 32'h00000000 /* 0xd4ac */;
                13612: data_o = 32'h00000000 /* 0xd4b0 */;
                13613: data_o = 32'h00000000 /* 0xd4b4 */;
                13614: data_o = 32'h00000000 /* 0xd4b8 */;
                13615: data_o = 32'h00000000 /* 0xd4bc */;
                13616: data_o = 32'h00000000 /* 0xd4c0 */;
                13617: data_o = 32'h00000000 /* 0xd4c4 */;
                13618: data_o = 32'h00000000 /* 0xd4c8 */;
                13619: data_o = 32'h00000000 /* 0xd4cc */;
                13620: data_o = 32'h00000000 /* 0xd4d0 */;
                13621: data_o = 32'h00000000 /* 0xd4d4 */;
                13622: data_o = 32'h00000000 /* 0xd4d8 */;
                13623: data_o = 32'h00000000 /* 0xd4dc */;
                13624: data_o = 32'h00000000 /* 0xd4e0 */;
                13625: data_o = 32'h00000000 /* 0xd4e4 */;
                13626: data_o = 32'h00000000 /* 0xd4e8 */;
                13627: data_o = 32'h00000000 /* 0xd4ec */;
                13628: data_o = 32'h00000000 /* 0xd4f0 */;
                13629: data_o = 32'h00000000 /* 0xd4f4 */;
                13630: data_o = 32'h00000000 /* 0xd4f8 */;
                13631: data_o = 32'h00000000 /* 0xd4fc */;
                13632: data_o = 32'h00000000 /* 0xd500 */;
                13633: data_o = 32'h00000000 /* 0xd504 */;
                13634: data_o = 32'h00000000 /* 0xd508 */;
                13635: data_o = 32'h00000000 /* 0xd50c */;
                13636: data_o = 32'h00000000 /* 0xd510 */;
                13637: data_o = 32'h00000000 /* 0xd514 */;
                13638: data_o = 32'h00000000 /* 0xd518 */;
                13639: data_o = 32'h00000000 /* 0xd51c */;
                13640: data_o = 32'h00000000 /* 0xd520 */;
                13641: data_o = 32'h00000000 /* 0xd524 */;
                13642: data_o = 32'h00000000 /* 0xd528 */;
                13643: data_o = 32'h00000000 /* 0xd52c */;
                13644: data_o = 32'h00000000 /* 0xd530 */;
                13645: data_o = 32'h00000000 /* 0xd534 */;
                13646: data_o = 32'h00000000 /* 0xd538 */;
                13647: data_o = 32'h00000000 /* 0xd53c */;
                13648: data_o = 32'h00000000 /* 0xd540 */;
                13649: data_o = 32'h00000000 /* 0xd544 */;
                13650: data_o = 32'h00000000 /* 0xd548 */;
                13651: data_o = 32'h00000000 /* 0xd54c */;
                13652: data_o = 32'h00000000 /* 0xd550 */;
                13653: data_o = 32'h00000000 /* 0xd554 */;
                13654: data_o = 32'h00000000 /* 0xd558 */;
                13655: data_o = 32'h00000000 /* 0xd55c */;
                13656: data_o = 32'h00000000 /* 0xd560 */;
                13657: data_o = 32'h00000000 /* 0xd564 */;
                13658: data_o = 32'h00000000 /* 0xd568 */;
                13659: data_o = 32'h00000000 /* 0xd56c */;
                13660: data_o = 32'h00000000 /* 0xd570 */;
                13661: data_o = 32'h00000000 /* 0xd574 */;
                13662: data_o = 32'h00000000 /* 0xd578 */;
                13663: data_o = 32'h00000000 /* 0xd57c */;
                13664: data_o = 32'h00000000 /* 0xd580 */;
                13665: data_o = 32'h00000000 /* 0xd584 */;
                13666: data_o = 32'h00000000 /* 0xd588 */;
                13667: data_o = 32'h00000000 /* 0xd58c */;
                13668: data_o = 32'h00000000 /* 0xd590 */;
                13669: data_o = 32'h00000000 /* 0xd594 */;
                13670: data_o = 32'h00000000 /* 0xd598 */;
                13671: data_o = 32'h00000000 /* 0xd59c */;
                13672: data_o = 32'h00000000 /* 0xd5a0 */;
                13673: data_o = 32'h00000000 /* 0xd5a4 */;
                13674: data_o = 32'h00000000 /* 0xd5a8 */;
                13675: data_o = 32'h00000000 /* 0xd5ac */;
                13676: data_o = 32'h00000000 /* 0xd5b0 */;
                13677: data_o = 32'h00000000 /* 0xd5b4 */;
                13678: data_o = 32'h00000000 /* 0xd5b8 */;
                13679: data_o = 32'h00000000 /* 0xd5bc */;
                13680: data_o = 32'h00000000 /* 0xd5c0 */;
                13681: data_o = 32'h00000000 /* 0xd5c4 */;
                13682: data_o = 32'h00000000 /* 0xd5c8 */;
                13683: data_o = 32'h00000000 /* 0xd5cc */;
                13684: data_o = 32'h00000000 /* 0xd5d0 */;
                13685: data_o = 32'h00000000 /* 0xd5d4 */;
                13686: data_o = 32'h00000000 /* 0xd5d8 */;
                13687: data_o = 32'h00000000 /* 0xd5dc */;
                13688: data_o = 32'h00000000 /* 0xd5e0 */;
                13689: data_o = 32'h00000000 /* 0xd5e4 */;
                13690: data_o = 32'h00000000 /* 0xd5e8 */;
                13691: data_o = 32'h00000000 /* 0xd5ec */;
                13692: data_o = 32'h00000000 /* 0xd5f0 */;
                13693: data_o = 32'h00000000 /* 0xd5f4 */;
                13694: data_o = 32'h00000000 /* 0xd5f8 */;
                13695: data_o = 32'h00000000 /* 0xd5fc */;
                13696: data_o = 32'h00000000 /* 0xd600 */;
                13697: data_o = 32'h00000000 /* 0xd604 */;
                13698: data_o = 32'h00000000 /* 0xd608 */;
                13699: data_o = 32'h00000000 /* 0xd60c */;
                13700: data_o = 32'h00000000 /* 0xd610 */;
                13701: data_o = 32'h00000000 /* 0xd614 */;
                13702: data_o = 32'h00000000 /* 0xd618 */;
                13703: data_o = 32'h00000000 /* 0xd61c */;
                13704: data_o = 32'h00000000 /* 0xd620 */;
                13705: data_o = 32'h00000000 /* 0xd624 */;
                13706: data_o = 32'h00000000 /* 0xd628 */;
                13707: data_o = 32'h00000000 /* 0xd62c */;
                13708: data_o = 32'h00000000 /* 0xd630 */;
                13709: data_o = 32'h00000000 /* 0xd634 */;
                13710: data_o = 32'h00000000 /* 0xd638 */;
                13711: data_o = 32'h00000000 /* 0xd63c */;
                13712: data_o = 32'h00000000 /* 0xd640 */;
                13713: data_o = 32'h00000000 /* 0xd644 */;
                13714: data_o = 32'h00000000 /* 0xd648 */;
                13715: data_o = 32'h00000000 /* 0xd64c */;
                13716: data_o = 32'h00000000 /* 0xd650 */;
                13717: data_o = 32'h00000000 /* 0xd654 */;
                13718: data_o = 32'h00000000 /* 0xd658 */;
                13719: data_o = 32'h00000000 /* 0xd65c */;
                13720: data_o = 32'h00000000 /* 0xd660 */;
                13721: data_o = 32'h00000000 /* 0xd664 */;
                13722: data_o = 32'h00000000 /* 0xd668 */;
                13723: data_o = 32'h00000000 /* 0xd66c */;
                13724: data_o = 32'h00000000 /* 0xd670 */;
                13725: data_o = 32'h00000000 /* 0xd674 */;
                13726: data_o = 32'h00000000 /* 0xd678 */;
                13727: data_o = 32'h00000000 /* 0xd67c */;
                13728: data_o = 32'h00000000 /* 0xd680 */;
                13729: data_o = 32'h00000000 /* 0xd684 */;
                13730: data_o = 32'h00000000 /* 0xd688 */;
                13731: data_o = 32'h00000000 /* 0xd68c */;
                13732: data_o = 32'h00000000 /* 0xd690 */;
                13733: data_o = 32'h00000000 /* 0xd694 */;
                13734: data_o = 32'h00000000 /* 0xd698 */;
                13735: data_o = 32'h00000000 /* 0xd69c */;
                13736: data_o = 32'h00000000 /* 0xd6a0 */;
                13737: data_o = 32'h00000000 /* 0xd6a4 */;
                13738: data_o = 32'h00000000 /* 0xd6a8 */;
                13739: data_o = 32'h00000000 /* 0xd6ac */;
                13740: data_o = 32'h00000000 /* 0xd6b0 */;
                13741: data_o = 32'h00000000 /* 0xd6b4 */;
                13742: data_o = 32'h00000000 /* 0xd6b8 */;
                13743: data_o = 32'h00000000 /* 0xd6bc */;
                13744: data_o = 32'h00000000 /* 0xd6c0 */;
                13745: data_o = 32'h00000000 /* 0xd6c4 */;
                13746: data_o = 32'h00000000 /* 0xd6c8 */;
                13747: data_o = 32'h00000000 /* 0xd6cc */;
                13748: data_o = 32'h00000000 /* 0xd6d0 */;
                13749: data_o = 32'h00000000 /* 0xd6d4 */;
                13750: data_o = 32'h00000000 /* 0xd6d8 */;
                13751: data_o = 32'h00000000 /* 0xd6dc */;
                13752: data_o = 32'h00000000 /* 0xd6e0 */;
                13753: data_o = 32'h00000000 /* 0xd6e4 */;
                13754: data_o = 32'h00000000 /* 0xd6e8 */;
                13755: data_o = 32'h00000000 /* 0xd6ec */;
                13756: data_o = 32'h00000000 /* 0xd6f0 */;
                13757: data_o = 32'h00000000 /* 0xd6f4 */;
                13758: data_o = 32'h00000000 /* 0xd6f8 */;
                13759: data_o = 32'h00000000 /* 0xd6fc */;
                13760: data_o = 32'h00000000 /* 0xd700 */;
                13761: data_o = 32'h00000000 /* 0xd704 */;
                13762: data_o = 32'h00000000 /* 0xd708 */;
                13763: data_o = 32'h00000000 /* 0xd70c */;
                13764: data_o = 32'h00000000 /* 0xd710 */;
                13765: data_o = 32'h00000000 /* 0xd714 */;
                13766: data_o = 32'h00000000 /* 0xd718 */;
                13767: data_o = 32'h00000000 /* 0xd71c */;
                13768: data_o = 32'h00000000 /* 0xd720 */;
                13769: data_o = 32'h00000000 /* 0xd724 */;
                13770: data_o = 32'h00000000 /* 0xd728 */;
                13771: data_o = 32'h00000000 /* 0xd72c */;
                13772: data_o = 32'h00000000 /* 0xd730 */;
                13773: data_o = 32'h00000000 /* 0xd734 */;
                13774: data_o = 32'h00000000 /* 0xd738 */;
                13775: data_o = 32'h00000000 /* 0xd73c */;
                13776: data_o = 32'h00000000 /* 0xd740 */;
                13777: data_o = 32'h00000000 /* 0xd744 */;
                13778: data_o = 32'h00000000 /* 0xd748 */;
                13779: data_o = 32'h00000000 /* 0xd74c */;
                13780: data_o = 32'h00000000 /* 0xd750 */;
                13781: data_o = 32'h00000000 /* 0xd754 */;
                13782: data_o = 32'h00000000 /* 0xd758 */;
                13783: data_o = 32'h00000000 /* 0xd75c */;
                13784: data_o = 32'h00000000 /* 0xd760 */;
                13785: data_o = 32'h00000000 /* 0xd764 */;
                13786: data_o = 32'h00000000 /* 0xd768 */;
                13787: data_o = 32'h00000000 /* 0xd76c */;
                13788: data_o = 32'h00000000 /* 0xd770 */;
                13789: data_o = 32'h00000000 /* 0xd774 */;
                13790: data_o = 32'h00000000 /* 0xd778 */;
                13791: data_o = 32'h00000000 /* 0xd77c */;
                13792: data_o = 32'h00000000 /* 0xd780 */;
                13793: data_o = 32'h00000000 /* 0xd784 */;
                13794: data_o = 32'h00000000 /* 0xd788 */;
                13795: data_o = 32'h00000000 /* 0xd78c */;
                13796: data_o = 32'h00000000 /* 0xd790 */;
                13797: data_o = 32'h00000000 /* 0xd794 */;
                13798: data_o = 32'h00000000 /* 0xd798 */;
                13799: data_o = 32'h00000000 /* 0xd79c */;
                13800: data_o = 32'h00000000 /* 0xd7a0 */;
                13801: data_o = 32'h00000000 /* 0xd7a4 */;
                13802: data_o = 32'h00000000 /* 0xd7a8 */;
                13803: data_o = 32'h00000000 /* 0xd7ac */;
                13804: data_o = 32'h00000000 /* 0xd7b0 */;
                13805: data_o = 32'h00000000 /* 0xd7b4 */;
                13806: data_o = 32'h00000000 /* 0xd7b8 */;
                13807: data_o = 32'h00000000 /* 0xd7bc */;
                13808: data_o = 32'h00000000 /* 0xd7c0 */;
                13809: data_o = 32'h00000000 /* 0xd7c4 */;
                13810: data_o = 32'h00000000 /* 0xd7c8 */;
                13811: data_o = 32'h00000000 /* 0xd7cc */;
                13812: data_o = 32'h00000000 /* 0xd7d0 */;
                13813: data_o = 32'h00000000 /* 0xd7d4 */;
                13814: data_o = 32'h00000000 /* 0xd7d8 */;
                13815: data_o = 32'h00000000 /* 0xd7dc */;
                13816: data_o = 32'h00000000 /* 0xd7e0 */;
                13817: data_o = 32'h00000000 /* 0xd7e4 */;
                13818: data_o = 32'h00000000 /* 0xd7e8 */;
                13819: data_o = 32'h00000000 /* 0xd7ec */;
                13820: data_o = 32'h00000000 /* 0xd7f0 */;
                13821: data_o = 32'h00000000 /* 0xd7f4 */;
                13822: data_o = 32'h00000000 /* 0xd7f8 */;
                13823: data_o = 32'h00000000 /* 0xd7fc */;
                13824: data_o = 32'h00000000 /* 0xd800 */;
                13825: data_o = 32'h00000000 /* 0xd804 */;
                13826: data_o = 32'h00000000 /* 0xd808 */;
                13827: data_o = 32'h00000000 /* 0xd80c */;
                13828: data_o = 32'h00000000 /* 0xd810 */;
                13829: data_o = 32'h00000000 /* 0xd814 */;
                13830: data_o = 32'h00000000 /* 0xd818 */;
                13831: data_o = 32'h00000000 /* 0xd81c */;
                13832: data_o = 32'h00000000 /* 0xd820 */;
                13833: data_o = 32'h00000000 /* 0xd824 */;
                13834: data_o = 32'h00000000 /* 0xd828 */;
                13835: data_o = 32'h00000000 /* 0xd82c */;
                13836: data_o = 32'h00000000 /* 0xd830 */;
                13837: data_o = 32'h00000000 /* 0xd834 */;
                13838: data_o = 32'h00000000 /* 0xd838 */;
                13839: data_o = 32'h00000000 /* 0xd83c */;
                13840: data_o = 32'h00000000 /* 0xd840 */;
                13841: data_o = 32'h00000000 /* 0xd844 */;
                13842: data_o = 32'h00000000 /* 0xd848 */;
                13843: data_o = 32'h00000000 /* 0xd84c */;
                13844: data_o = 32'h00000000 /* 0xd850 */;
                13845: data_o = 32'h00000000 /* 0xd854 */;
                13846: data_o = 32'h00000000 /* 0xd858 */;
                13847: data_o = 32'h00000000 /* 0xd85c */;
                13848: data_o = 32'h00000000 /* 0xd860 */;
                13849: data_o = 32'h00000000 /* 0xd864 */;
                13850: data_o = 32'h00000000 /* 0xd868 */;
                13851: data_o = 32'h00000000 /* 0xd86c */;
                13852: data_o = 32'h00000000 /* 0xd870 */;
                13853: data_o = 32'h00000000 /* 0xd874 */;
                13854: data_o = 32'h00000000 /* 0xd878 */;
                13855: data_o = 32'h00000000 /* 0xd87c */;
                13856: data_o = 32'h00000000 /* 0xd880 */;
                13857: data_o = 32'h00000000 /* 0xd884 */;
                13858: data_o = 32'h00000000 /* 0xd888 */;
                13859: data_o = 32'h00000000 /* 0xd88c */;
                13860: data_o = 32'h00000000 /* 0xd890 */;
                13861: data_o = 32'h00000000 /* 0xd894 */;
                13862: data_o = 32'h00000000 /* 0xd898 */;
                13863: data_o = 32'h00000000 /* 0xd89c */;
                13864: data_o = 32'h00000000 /* 0xd8a0 */;
                13865: data_o = 32'h00000000 /* 0xd8a4 */;
                13866: data_o = 32'h00000000 /* 0xd8a8 */;
                13867: data_o = 32'h00000000 /* 0xd8ac */;
                13868: data_o = 32'h00000000 /* 0xd8b0 */;
                13869: data_o = 32'h00000000 /* 0xd8b4 */;
                13870: data_o = 32'h00000000 /* 0xd8b8 */;
                13871: data_o = 32'h00000000 /* 0xd8bc */;
                13872: data_o = 32'h00000000 /* 0xd8c0 */;
                13873: data_o = 32'h00000000 /* 0xd8c4 */;
                13874: data_o = 32'h00000000 /* 0xd8c8 */;
                13875: data_o = 32'h00000000 /* 0xd8cc */;
                13876: data_o = 32'h00000000 /* 0xd8d0 */;
                13877: data_o = 32'h00000000 /* 0xd8d4 */;
                13878: data_o = 32'h00000000 /* 0xd8d8 */;
                13879: data_o = 32'h00000000 /* 0xd8dc */;
                13880: data_o = 32'h00000000 /* 0xd8e0 */;
                13881: data_o = 32'h00000000 /* 0xd8e4 */;
                13882: data_o = 32'h00000000 /* 0xd8e8 */;
                13883: data_o = 32'h00000000 /* 0xd8ec */;
                13884: data_o = 32'h00000000 /* 0xd8f0 */;
                13885: data_o = 32'h00000000 /* 0xd8f4 */;
                13886: data_o = 32'h00000000 /* 0xd8f8 */;
                13887: data_o = 32'h00000000 /* 0xd8fc */;
                13888: data_o = 32'h00000000 /* 0xd900 */;
                13889: data_o = 32'h00000000 /* 0xd904 */;
                13890: data_o = 32'h00000000 /* 0xd908 */;
                13891: data_o = 32'h00000000 /* 0xd90c */;
                13892: data_o = 32'h00000000 /* 0xd910 */;
                13893: data_o = 32'h00000000 /* 0xd914 */;
                13894: data_o = 32'h00000000 /* 0xd918 */;
                13895: data_o = 32'h00000000 /* 0xd91c */;
                13896: data_o = 32'h00000000 /* 0xd920 */;
                13897: data_o = 32'h00000000 /* 0xd924 */;
                13898: data_o = 32'h00000000 /* 0xd928 */;
                13899: data_o = 32'h00000000 /* 0xd92c */;
                13900: data_o = 32'h00000000 /* 0xd930 */;
                13901: data_o = 32'h00000000 /* 0xd934 */;
                13902: data_o = 32'h00000000 /* 0xd938 */;
                13903: data_o = 32'h00000000 /* 0xd93c */;
                13904: data_o = 32'h00000000 /* 0xd940 */;
                13905: data_o = 32'h00000000 /* 0xd944 */;
                13906: data_o = 32'h00000000 /* 0xd948 */;
                13907: data_o = 32'h00000000 /* 0xd94c */;
                13908: data_o = 32'h00000000 /* 0xd950 */;
                13909: data_o = 32'h00000000 /* 0xd954 */;
                13910: data_o = 32'h00000000 /* 0xd958 */;
                13911: data_o = 32'h00000000 /* 0xd95c */;
                13912: data_o = 32'h00000000 /* 0xd960 */;
                13913: data_o = 32'h00000000 /* 0xd964 */;
                13914: data_o = 32'h00000000 /* 0xd968 */;
                13915: data_o = 32'h00000000 /* 0xd96c */;
                13916: data_o = 32'h00000000 /* 0xd970 */;
                13917: data_o = 32'h00000000 /* 0xd974 */;
                13918: data_o = 32'h00000000 /* 0xd978 */;
                13919: data_o = 32'h00000000 /* 0xd97c */;
                13920: data_o = 32'h00000000 /* 0xd980 */;
                13921: data_o = 32'h00000000 /* 0xd984 */;
                13922: data_o = 32'h00000000 /* 0xd988 */;
                13923: data_o = 32'h00000000 /* 0xd98c */;
                13924: data_o = 32'h00000000 /* 0xd990 */;
                13925: data_o = 32'h00000000 /* 0xd994 */;
                13926: data_o = 32'h00000000 /* 0xd998 */;
                13927: data_o = 32'h00000000 /* 0xd99c */;
                13928: data_o = 32'h00000000 /* 0xd9a0 */;
                13929: data_o = 32'h00000000 /* 0xd9a4 */;
                13930: data_o = 32'h00000000 /* 0xd9a8 */;
                13931: data_o = 32'h00000000 /* 0xd9ac */;
                13932: data_o = 32'h00000000 /* 0xd9b0 */;
                13933: data_o = 32'h00000000 /* 0xd9b4 */;
                13934: data_o = 32'h00000000 /* 0xd9b8 */;
                13935: data_o = 32'h00000000 /* 0xd9bc */;
                13936: data_o = 32'h00000000 /* 0xd9c0 */;
                13937: data_o = 32'h00000000 /* 0xd9c4 */;
                13938: data_o = 32'h00000000 /* 0xd9c8 */;
                13939: data_o = 32'h00000000 /* 0xd9cc */;
                13940: data_o = 32'h00000000 /* 0xd9d0 */;
                13941: data_o = 32'h00000000 /* 0xd9d4 */;
                13942: data_o = 32'h00000000 /* 0xd9d8 */;
                13943: data_o = 32'h00000000 /* 0xd9dc */;
                13944: data_o = 32'h00000000 /* 0xd9e0 */;
                13945: data_o = 32'h00000000 /* 0xd9e4 */;
                13946: data_o = 32'h00000000 /* 0xd9e8 */;
                13947: data_o = 32'h00000000 /* 0xd9ec */;
                13948: data_o = 32'h00000000 /* 0xd9f0 */;
                13949: data_o = 32'h00000000 /* 0xd9f4 */;
                13950: data_o = 32'h00000000 /* 0xd9f8 */;
                13951: data_o = 32'h00000000 /* 0xd9fc */;
                13952: data_o = 32'h00000000 /* 0xda00 */;
                13953: data_o = 32'h00000000 /* 0xda04 */;
                13954: data_o = 32'h00000000 /* 0xda08 */;
                13955: data_o = 32'h00000000 /* 0xda0c */;
                13956: data_o = 32'h00000000 /* 0xda10 */;
                13957: data_o = 32'h00000000 /* 0xda14 */;
                13958: data_o = 32'h00000000 /* 0xda18 */;
                13959: data_o = 32'h00000000 /* 0xda1c */;
                13960: data_o = 32'h00000000 /* 0xda20 */;
                13961: data_o = 32'h00000000 /* 0xda24 */;
                13962: data_o = 32'h00000000 /* 0xda28 */;
                13963: data_o = 32'h00000000 /* 0xda2c */;
                13964: data_o = 32'h00000000 /* 0xda30 */;
                13965: data_o = 32'h00000000 /* 0xda34 */;
                13966: data_o = 32'h00000000 /* 0xda38 */;
                13967: data_o = 32'h00000000 /* 0xda3c */;
                13968: data_o = 32'h00000000 /* 0xda40 */;
                13969: data_o = 32'h00000000 /* 0xda44 */;
                13970: data_o = 32'h00000000 /* 0xda48 */;
                13971: data_o = 32'h00000000 /* 0xda4c */;
                13972: data_o = 32'h00000000 /* 0xda50 */;
                13973: data_o = 32'h00000000 /* 0xda54 */;
                13974: data_o = 32'h00000000 /* 0xda58 */;
                13975: data_o = 32'h00000000 /* 0xda5c */;
                13976: data_o = 32'h00000000 /* 0xda60 */;
                13977: data_o = 32'h00000000 /* 0xda64 */;
                13978: data_o = 32'h00000000 /* 0xda68 */;
                13979: data_o = 32'h00000000 /* 0xda6c */;
                13980: data_o = 32'h00000000 /* 0xda70 */;
                13981: data_o = 32'h00000000 /* 0xda74 */;
                13982: data_o = 32'h00000000 /* 0xda78 */;
                13983: data_o = 32'h00000000 /* 0xda7c */;
                13984: data_o = 32'h00000000 /* 0xda80 */;
                13985: data_o = 32'h00000000 /* 0xda84 */;
                13986: data_o = 32'h00000000 /* 0xda88 */;
                13987: data_o = 32'h00000000 /* 0xda8c */;
                13988: data_o = 32'h00000000 /* 0xda90 */;
                13989: data_o = 32'h00000000 /* 0xda94 */;
                13990: data_o = 32'h00000000 /* 0xda98 */;
                13991: data_o = 32'h00000000 /* 0xda9c */;
                13992: data_o = 32'h00000000 /* 0xdaa0 */;
                13993: data_o = 32'h00000000 /* 0xdaa4 */;
                13994: data_o = 32'h00000000 /* 0xdaa8 */;
                13995: data_o = 32'h00000000 /* 0xdaac */;
                13996: data_o = 32'h00000000 /* 0xdab0 */;
                13997: data_o = 32'h00000000 /* 0xdab4 */;
                13998: data_o = 32'h00000000 /* 0xdab8 */;
                13999: data_o = 32'h00000000 /* 0xdabc */;
                14000: data_o = 32'h00000000 /* 0xdac0 */;
                14001: data_o = 32'h00000000 /* 0xdac4 */;
                14002: data_o = 32'h00000000 /* 0xdac8 */;
                14003: data_o = 32'h00000000 /* 0xdacc */;
                14004: data_o = 32'h00000000 /* 0xdad0 */;
                14005: data_o = 32'h00000000 /* 0xdad4 */;
                14006: data_o = 32'h00000000 /* 0xdad8 */;
                14007: data_o = 32'h00000000 /* 0xdadc */;
                14008: data_o = 32'h00000000 /* 0xdae0 */;
                14009: data_o = 32'h00000000 /* 0xdae4 */;
                14010: data_o = 32'h00000000 /* 0xdae8 */;
                14011: data_o = 32'h00000000 /* 0xdaec */;
                14012: data_o = 32'h00000000 /* 0xdaf0 */;
                14013: data_o = 32'h00000000 /* 0xdaf4 */;
                14014: data_o = 32'h00000000 /* 0xdaf8 */;
                14015: data_o = 32'h00000000 /* 0xdafc */;
                14016: data_o = 32'h00000000 /* 0xdb00 */;
                14017: data_o = 32'h00000000 /* 0xdb04 */;
                14018: data_o = 32'h00000000 /* 0xdb08 */;
                14019: data_o = 32'h00000000 /* 0xdb0c */;
                14020: data_o = 32'h00000000 /* 0xdb10 */;
                14021: data_o = 32'h00000000 /* 0xdb14 */;
                14022: data_o = 32'h00000000 /* 0xdb18 */;
                14023: data_o = 32'h00000000 /* 0xdb1c */;
                14024: data_o = 32'h00000000 /* 0xdb20 */;
                14025: data_o = 32'h00000000 /* 0xdb24 */;
                14026: data_o = 32'h00000000 /* 0xdb28 */;
                14027: data_o = 32'h00000000 /* 0xdb2c */;
                14028: data_o = 32'h00000000 /* 0xdb30 */;
                14029: data_o = 32'h00000000 /* 0xdb34 */;
                14030: data_o = 32'h00000000 /* 0xdb38 */;
                14031: data_o = 32'h00000000 /* 0xdb3c */;
                14032: data_o = 32'h00000000 /* 0xdb40 */;
                14033: data_o = 32'h00000000 /* 0xdb44 */;
                14034: data_o = 32'h00000000 /* 0xdb48 */;
                14035: data_o = 32'h00000000 /* 0xdb4c */;
                14036: data_o = 32'h00000000 /* 0xdb50 */;
                14037: data_o = 32'h00000000 /* 0xdb54 */;
                14038: data_o = 32'h00000000 /* 0xdb58 */;
                14039: data_o = 32'h00000000 /* 0xdb5c */;
                14040: data_o = 32'h00000000 /* 0xdb60 */;
                14041: data_o = 32'h00000000 /* 0xdb64 */;
                14042: data_o = 32'h00000000 /* 0xdb68 */;
                14043: data_o = 32'h00000000 /* 0xdb6c */;
                14044: data_o = 32'h00000000 /* 0xdb70 */;
                14045: data_o = 32'h00000000 /* 0xdb74 */;
                14046: data_o = 32'h00000000 /* 0xdb78 */;
                14047: data_o = 32'h00000000 /* 0xdb7c */;
                14048: data_o = 32'h00000000 /* 0xdb80 */;
                14049: data_o = 32'h00000000 /* 0xdb84 */;
                14050: data_o = 32'h00000000 /* 0xdb88 */;
                14051: data_o = 32'h00000000 /* 0xdb8c */;
                14052: data_o = 32'h00000000 /* 0xdb90 */;
                14053: data_o = 32'h00000000 /* 0xdb94 */;
                14054: data_o = 32'h00000000 /* 0xdb98 */;
                14055: data_o = 32'h00000000 /* 0xdb9c */;
                14056: data_o = 32'h00000000 /* 0xdba0 */;
                14057: data_o = 32'h00000000 /* 0xdba4 */;
                14058: data_o = 32'h00000000 /* 0xdba8 */;
                14059: data_o = 32'h00000000 /* 0xdbac */;
                14060: data_o = 32'h00000000 /* 0xdbb0 */;
                14061: data_o = 32'h00000000 /* 0xdbb4 */;
                14062: data_o = 32'h00000000 /* 0xdbb8 */;
                14063: data_o = 32'h00000000 /* 0xdbbc */;
                14064: data_o = 32'h00000000 /* 0xdbc0 */;
                14065: data_o = 32'h00000000 /* 0xdbc4 */;
                14066: data_o = 32'h00000000 /* 0xdbc8 */;
                14067: data_o = 32'h00000000 /* 0xdbcc */;
                14068: data_o = 32'h00000000 /* 0xdbd0 */;
                14069: data_o = 32'h00000000 /* 0xdbd4 */;
                14070: data_o = 32'h00000000 /* 0xdbd8 */;
                14071: data_o = 32'h00000000 /* 0xdbdc */;
                14072: data_o = 32'h00000000 /* 0xdbe0 */;
                14073: data_o = 32'h00000000 /* 0xdbe4 */;
                14074: data_o = 32'h00000000 /* 0xdbe8 */;
                14075: data_o = 32'h00000000 /* 0xdbec */;
                14076: data_o = 32'h00000000 /* 0xdbf0 */;
                14077: data_o = 32'h00000000 /* 0xdbf4 */;
                14078: data_o = 32'h00000000 /* 0xdbf8 */;
                14079: data_o = 32'h00000000 /* 0xdbfc */;
                14080: data_o = 32'h00000000 /* 0xdc00 */;
                14081: data_o = 32'h00000000 /* 0xdc04 */;
                14082: data_o = 32'h00000000 /* 0xdc08 */;
                14083: data_o = 32'h00000000 /* 0xdc0c */;
                14084: data_o = 32'h00000000 /* 0xdc10 */;
                14085: data_o = 32'h00000000 /* 0xdc14 */;
                14086: data_o = 32'h00000000 /* 0xdc18 */;
                14087: data_o = 32'h00000000 /* 0xdc1c */;
                14088: data_o = 32'h00000000 /* 0xdc20 */;
                14089: data_o = 32'h00000000 /* 0xdc24 */;
                14090: data_o = 32'h00000000 /* 0xdc28 */;
                14091: data_o = 32'h00000000 /* 0xdc2c */;
                14092: data_o = 32'h00000000 /* 0xdc30 */;
                14093: data_o = 32'h00000000 /* 0xdc34 */;
                14094: data_o = 32'h00000000 /* 0xdc38 */;
                14095: data_o = 32'h00000000 /* 0xdc3c */;
                14096: data_o = 32'h00000000 /* 0xdc40 */;
                14097: data_o = 32'h00000000 /* 0xdc44 */;
                14098: data_o = 32'h00000000 /* 0xdc48 */;
                14099: data_o = 32'h00000000 /* 0xdc4c */;
                14100: data_o = 32'h00000000 /* 0xdc50 */;
                14101: data_o = 32'h00000000 /* 0xdc54 */;
                14102: data_o = 32'h00000000 /* 0xdc58 */;
                14103: data_o = 32'h00000000 /* 0xdc5c */;
                14104: data_o = 32'h00000000 /* 0xdc60 */;
                14105: data_o = 32'h00000000 /* 0xdc64 */;
                14106: data_o = 32'h00000000 /* 0xdc68 */;
                14107: data_o = 32'h00000000 /* 0xdc6c */;
                14108: data_o = 32'h00000000 /* 0xdc70 */;
                14109: data_o = 32'h00000000 /* 0xdc74 */;
                14110: data_o = 32'h00000000 /* 0xdc78 */;
                14111: data_o = 32'h00000000 /* 0xdc7c */;
                14112: data_o = 32'h00000000 /* 0xdc80 */;
                14113: data_o = 32'h00000000 /* 0xdc84 */;
                14114: data_o = 32'h00000000 /* 0xdc88 */;
                14115: data_o = 32'h00000000 /* 0xdc8c */;
                14116: data_o = 32'h00000000 /* 0xdc90 */;
                14117: data_o = 32'h00000000 /* 0xdc94 */;
                14118: data_o = 32'h00000000 /* 0xdc98 */;
                14119: data_o = 32'h00000000 /* 0xdc9c */;
                14120: data_o = 32'h00000000 /* 0xdca0 */;
                14121: data_o = 32'h00000000 /* 0xdca4 */;
                14122: data_o = 32'h00000000 /* 0xdca8 */;
                14123: data_o = 32'h00000000 /* 0xdcac */;
                14124: data_o = 32'h00000000 /* 0xdcb0 */;
                14125: data_o = 32'h00000000 /* 0xdcb4 */;
                14126: data_o = 32'h00000000 /* 0xdcb8 */;
                14127: data_o = 32'h00000000 /* 0xdcbc */;
                14128: data_o = 32'h00000000 /* 0xdcc0 */;
                14129: data_o = 32'h00000000 /* 0xdcc4 */;
                14130: data_o = 32'h00000000 /* 0xdcc8 */;
                14131: data_o = 32'h00000000 /* 0xdccc */;
                14132: data_o = 32'h00000000 /* 0xdcd0 */;
                14133: data_o = 32'h00000000 /* 0xdcd4 */;
                14134: data_o = 32'h00000000 /* 0xdcd8 */;
                14135: data_o = 32'h00000000 /* 0xdcdc */;
                14136: data_o = 32'h00000000 /* 0xdce0 */;
                14137: data_o = 32'h00000000 /* 0xdce4 */;
                14138: data_o = 32'h00000000 /* 0xdce8 */;
                14139: data_o = 32'h00000000 /* 0xdcec */;
                14140: data_o = 32'h00000000 /* 0xdcf0 */;
                14141: data_o = 32'h00000000 /* 0xdcf4 */;
                14142: data_o = 32'h00000000 /* 0xdcf8 */;
                14143: data_o = 32'h00000000 /* 0xdcfc */;
                14144: data_o = 32'h00000000 /* 0xdd00 */;
                14145: data_o = 32'h00000000 /* 0xdd04 */;
                14146: data_o = 32'h00000000 /* 0xdd08 */;
                14147: data_o = 32'h00000000 /* 0xdd0c */;
                14148: data_o = 32'h00000000 /* 0xdd10 */;
                14149: data_o = 32'h00000000 /* 0xdd14 */;
                14150: data_o = 32'h00000000 /* 0xdd18 */;
                14151: data_o = 32'h00000000 /* 0xdd1c */;
                14152: data_o = 32'h00000000 /* 0xdd20 */;
                14153: data_o = 32'h00000000 /* 0xdd24 */;
                14154: data_o = 32'h00000000 /* 0xdd28 */;
                14155: data_o = 32'h00000000 /* 0xdd2c */;
                14156: data_o = 32'h00000000 /* 0xdd30 */;
                14157: data_o = 32'h00000000 /* 0xdd34 */;
                14158: data_o = 32'h00000000 /* 0xdd38 */;
                14159: data_o = 32'h00000000 /* 0xdd3c */;
                14160: data_o = 32'h00000000 /* 0xdd40 */;
                14161: data_o = 32'h00000000 /* 0xdd44 */;
                14162: data_o = 32'h00000000 /* 0xdd48 */;
                14163: data_o = 32'h00000000 /* 0xdd4c */;
                14164: data_o = 32'h00000000 /* 0xdd50 */;
                14165: data_o = 32'h00000000 /* 0xdd54 */;
                14166: data_o = 32'h00000000 /* 0xdd58 */;
                14167: data_o = 32'h00000000 /* 0xdd5c */;
                14168: data_o = 32'h00000000 /* 0xdd60 */;
                14169: data_o = 32'h00000000 /* 0xdd64 */;
                14170: data_o = 32'h00000000 /* 0xdd68 */;
                14171: data_o = 32'h00000000 /* 0xdd6c */;
                14172: data_o = 32'h00000000 /* 0xdd70 */;
                14173: data_o = 32'h00000000 /* 0xdd74 */;
                14174: data_o = 32'h00000000 /* 0xdd78 */;
                14175: data_o = 32'h00000000 /* 0xdd7c */;
                14176: data_o = 32'h00000000 /* 0xdd80 */;
                14177: data_o = 32'h00000000 /* 0xdd84 */;
                14178: data_o = 32'h00000000 /* 0xdd88 */;
                14179: data_o = 32'h00000000 /* 0xdd8c */;
                14180: data_o = 32'h00000000 /* 0xdd90 */;
                14181: data_o = 32'h00000000 /* 0xdd94 */;
                14182: data_o = 32'h00000000 /* 0xdd98 */;
                14183: data_o = 32'h00000000 /* 0xdd9c */;
                14184: data_o = 32'h00000000 /* 0xdda0 */;
                14185: data_o = 32'h00000000 /* 0xdda4 */;
                14186: data_o = 32'h00000000 /* 0xdda8 */;
                14187: data_o = 32'h00000000 /* 0xddac */;
                14188: data_o = 32'h00000000 /* 0xddb0 */;
                14189: data_o = 32'h00000000 /* 0xddb4 */;
                14190: data_o = 32'h00000000 /* 0xddb8 */;
                14191: data_o = 32'h00000000 /* 0xddbc */;
                14192: data_o = 32'h00000000 /* 0xddc0 */;
                14193: data_o = 32'h00000000 /* 0xddc4 */;
                14194: data_o = 32'h00000000 /* 0xddc8 */;
                14195: data_o = 32'h00000000 /* 0xddcc */;
                14196: data_o = 32'h00000000 /* 0xddd0 */;
                14197: data_o = 32'h00000000 /* 0xddd4 */;
                14198: data_o = 32'h00000000 /* 0xddd8 */;
                14199: data_o = 32'h00000000 /* 0xdddc */;
                14200: data_o = 32'h00000000 /* 0xdde0 */;
                14201: data_o = 32'h00000000 /* 0xdde4 */;
                14202: data_o = 32'h00000000 /* 0xdde8 */;
                14203: data_o = 32'h00000000 /* 0xddec */;
                14204: data_o = 32'h00000000 /* 0xddf0 */;
                14205: data_o = 32'h00000000 /* 0xddf4 */;
                14206: data_o = 32'h00000000 /* 0xddf8 */;
                14207: data_o = 32'h00000000 /* 0xddfc */;
                14208: data_o = 32'h00000000 /* 0xde00 */;
                14209: data_o = 32'h00000000 /* 0xde04 */;
                14210: data_o = 32'h00000000 /* 0xde08 */;
                14211: data_o = 32'h00000000 /* 0xde0c */;
                14212: data_o = 32'h00000000 /* 0xde10 */;
                14213: data_o = 32'h00000000 /* 0xde14 */;
                14214: data_o = 32'h00000000 /* 0xde18 */;
                14215: data_o = 32'h00000000 /* 0xde1c */;
                14216: data_o = 32'h00000000 /* 0xde20 */;
                14217: data_o = 32'h00000000 /* 0xde24 */;
                14218: data_o = 32'h00000000 /* 0xde28 */;
                14219: data_o = 32'h00000000 /* 0xde2c */;
                14220: data_o = 32'h00000000 /* 0xde30 */;
                14221: data_o = 32'h00000000 /* 0xde34 */;
                14222: data_o = 32'h00000000 /* 0xde38 */;
                14223: data_o = 32'h00000000 /* 0xde3c */;
                14224: data_o = 32'h00000000 /* 0xde40 */;
                14225: data_o = 32'h00000000 /* 0xde44 */;
                14226: data_o = 32'h00000000 /* 0xde48 */;
                14227: data_o = 32'h00000000 /* 0xde4c */;
                14228: data_o = 32'h00000000 /* 0xde50 */;
                14229: data_o = 32'h00000000 /* 0xde54 */;
                14230: data_o = 32'h00000000 /* 0xde58 */;
                14231: data_o = 32'h00000000 /* 0xde5c */;
                14232: data_o = 32'h00000000 /* 0xde60 */;
                14233: data_o = 32'h00000000 /* 0xde64 */;
                14234: data_o = 32'h00000000 /* 0xde68 */;
                14235: data_o = 32'h00000000 /* 0xde6c */;
                14236: data_o = 32'h00000000 /* 0xde70 */;
                14237: data_o = 32'h00000000 /* 0xde74 */;
                14238: data_o = 32'h00000000 /* 0xde78 */;
                14239: data_o = 32'h00000000 /* 0xde7c */;
                14240: data_o = 32'h00000000 /* 0xde80 */;
                14241: data_o = 32'h00000000 /* 0xde84 */;
                14242: data_o = 32'h00000000 /* 0xde88 */;
                14243: data_o = 32'h00000000 /* 0xde8c */;
                14244: data_o = 32'h00000000 /* 0xde90 */;
                14245: data_o = 32'h00000000 /* 0xde94 */;
                14246: data_o = 32'h00000000 /* 0xde98 */;
                14247: data_o = 32'h00000000 /* 0xde9c */;
                14248: data_o = 32'h00000000 /* 0xdea0 */;
                14249: data_o = 32'h00000000 /* 0xdea4 */;
                14250: data_o = 32'h00000000 /* 0xdea8 */;
                14251: data_o = 32'h00000000 /* 0xdeac */;
                14252: data_o = 32'h00000000 /* 0xdeb0 */;
                14253: data_o = 32'h00000000 /* 0xdeb4 */;
                14254: data_o = 32'h00000000 /* 0xdeb8 */;
                14255: data_o = 32'h00000000 /* 0xdebc */;
                14256: data_o = 32'h00000000 /* 0xdec0 */;
                14257: data_o = 32'h00000000 /* 0xdec4 */;
                14258: data_o = 32'h00000000 /* 0xdec8 */;
                14259: data_o = 32'h00000000 /* 0xdecc */;
                14260: data_o = 32'h00000000 /* 0xded0 */;
                14261: data_o = 32'h00000000 /* 0xded4 */;
                14262: data_o = 32'h00000000 /* 0xded8 */;
                14263: data_o = 32'h00000000 /* 0xdedc */;
                14264: data_o = 32'h00000000 /* 0xdee0 */;
                14265: data_o = 32'h00000000 /* 0xdee4 */;
                14266: data_o = 32'h00000000 /* 0xdee8 */;
                14267: data_o = 32'h00000000 /* 0xdeec */;
                14268: data_o = 32'h00000000 /* 0xdef0 */;
                14269: data_o = 32'h00000000 /* 0xdef4 */;
                14270: data_o = 32'h00000000 /* 0xdef8 */;
                14271: data_o = 32'h00000000 /* 0xdefc */;
                14272: data_o = 32'h00000000 /* 0xdf00 */;
                14273: data_o = 32'h00000000 /* 0xdf04 */;
                14274: data_o = 32'h00000000 /* 0xdf08 */;
                14275: data_o = 32'h00000000 /* 0xdf0c */;
                14276: data_o = 32'h00000000 /* 0xdf10 */;
                14277: data_o = 32'h00000000 /* 0xdf14 */;
                14278: data_o = 32'h00000000 /* 0xdf18 */;
                14279: data_o = 32'h00000000 /* 0xdf1c */;
                14280: data_o = 32'h00000000 /* 0xdf20 */;
                14281: data_o = 32'h00000000 /* 0xdf24 */;
                14282: data_o = 32'h00000000 /* 0xdf28 */;
                14283: data_o = 32'h00000000 /* 0xdf2c */;
                14284: data_o = 32'h00000000 /* 0xdf30 */;
                14285: data_o = 32'h00000000 /* 0xdf34 */;
                14286: data_o = 32'h00000000 /* 0xdf38 */;
                14287: data_o = 32'h00000000 /* 0xdf3c */;
                14288: data_o = 32'h00000000 /* 0xdf40 */;
                14289: data_o = 32'h00000000 /* 0xdf44 */;
                14290: data_o = 32'h00000000 /* 0xdf48 */;
                14291: data_o = 32'h00000000 /* 0xdf4c */;
                14292: data_o = 32'h00000000 /* 0xdf50 */;
                14293: data_o = 32'h00000000 /* 0xdf54 */;
                14294: data_o = 32'h00000000 /* 0xdf58 */;
                14295: data_o = 32'h00000000 /* 0xdf5c */;
                14296: data_o = 32'h00000000 /* 0xdf60 */;
                14297: data_o = 32'h00000000 /* 0xdf64 */;
                14298: data_o = 32'h00000000 /* 0xdf68 */;
                14299: data_o = 32'h00000000 /* 0xdf6c */;
                14300: data_o = 32'h00000000 /* 0xdf70 */;
                14301: data_o = 32'h00000000 /* 0xdf74 */;
                14302: data_o = 32'h00000000 /* 0xdf78 */;
                14303: data_o = 32'h00000000 /* 0xdf7c */;
                14304: data_o = 32'h00000000 /* 0xdf80 */;
                14305: data_o = 32'h00000000 /* 0xdf84 */;
                14306: data_o = 32'h00000000 /* 0xdf88 */;
                14307: data_o = 32'h00000000 /* 0xdf8c */;
                14308: data_o = 32'h00000000 /* 0xdf90 */;
                14309: data_o = 32'h00000000 /* 0xdf94 */;
                14310: data_o = 32'h00000000 /* 0xdf98 */;
                14311: data_o = 32'h00000000 /* 0xdf9c */;
                14312: data_o = 32'h00000000 /* 0xdfa0 */;
                14313: data_o = 32'h00000000 /* 0xdfa4 */;
                14314: data_o = 32'h00000000 /* 0xdfa8 */;
                14315: data_o = 32'h00000000 /* 0xdfac */;
                14316: data_o = 32'h00000000 /* 0xdfb0 */;
                14317: data_o = 32'h00000000 /* 0xdfb4 */;
                14318: data_o = 32'h00000000 /* 0xdfb8 */;
                14319: data_o = 32'h00000000 /* 0xdfbc */;
                14320: data_o = 32'h00000000 /* 0xdfc0 */;
                14321: data_o = 32'h00000000 /* 0xdfc4 */;
                14322: data_o = 32'h00000000 /* 0xdfc8 */;
                14323: data_o = 32'h00000000 /* 0xdfcc */;
                14324: data_o = 32'h00000000 /* 0xdfd0 */;
                14325: data_o = 32'h00000000 /* 0xdfd4 */;
                14326: data_o = 32'h00000000 /* 0xdfd8 */;
                14327: data_o = 32'h00000000 /* 0xdfdc */;
                14328: data_o = 32'h00000000 /* 0xdfe0 */;
                14329: data_o = 32'h00000000 /* 0xdfe4 */;
                14330: data_o = 32'h00000000 /* 0xdfe8 */;
                14331: data_o = 32'h00000000 /* 0xdfec */;
                14332: data_o = 32'h00000000 /* 0xdff0 */;
                14333: data_o = 32'h00000000 /* 0xdff4 */;
                14334: data_o = 32'h00000000 /* 0xdff8 */;
                14335: data_o = 32'h00000000 /* 0xdffc */;
                14336: data_o = 32'h00000000 /* 0xe000 */;
                14337: data_o = 32'h00000000 /* 0xe004 */;
                14338: data_o = 32'h00000000 /* 0xe008 */;
                14339: data_o = 32'h00000000 /* 0xe00c */;
                14340: data_o = 32'h00000000 /* 0xe010 */;
                14341: data_o = 32'h00000000 /* 0xe014 */;
                14342: data_o = 32'h00000000 /* 0xe018 */;
                14343: data_o = 32'h00000000 /* 0xe01c */;
                14344: data_o = 32'h00000000 /* 0xe020 */;
                14345: data_o = 32'h00000000 /* 0xe024 */;
                14346: data_o = 32'h00000000 /* 0xe028 */;
                14347: data_o = 32'h00000000 /* 0xe02c */;
                14348: data_o = 32'h00000000 /* 0xe030 */;
                14349: data_o = 32'h00000000 /* 0xe034 */;
                14350: data_o = 32'h00000000 /* 0xe038 */;
                14351: data_o = 32'h00000000 /* 0xe03c */;
                14352: data_o = 32'h00000000 /* 0xe040 */;
                14353: data_o = 32'h00000000 /* 0xe044 */;
                14354: data_o = 32'h00000000 /* 0xe048 */;
                14355: data_o = 32'h00000000 /* 0xe04c */;
                14356: data_o = 32'h00000000 /* 0xe050 */;
                14357: data_o = 32'h00000000 /* 0xe054 */;
                14358: data_o = 32'h00000000 /* 0xe058 */;
                14359: data_o = 32'h00000000 /* 0xe05c */;
                14360: data_o = 32'h00000000 /* 0xe060 */;
                14361: data_o = 32'h00000000 /* 0xe064 */;
                14362: data_o = 32'h00000000 /* 0xe068 */;
                14363: data_o = 32'h00000000 /* 0xe06c */;
                14364: data_o = 32'h00000000 /* 0xe070 */;
                14365: data_o = 32'h00000000 /* 0xe074 */;
                14366: data_o = 32'h00000000 /* 0xe078 */;
                14367: data_o = 32'h00000000 /* 0xe07c */;
                14368: data_o = 32'h00000000 /* 0xe080 */;
                14369: data_o = 32'h00000000 /* 0xe084 */;
                14370: data_o = 32'h00000000 /* 0xe088 */;
                14371: data_o = 32'h00000000 /* 0xe08c */;
                14372: data_o = 32'h00000000 /* 0xe090 */;
                14373: data_o = 32'h00000000 /* 0xe094 */;
                14374: data_o = 32'h00000000 /* 0xe098 */;
                14375: data_o = 32'h00000000 /* 0xe09c */;
                14376: data_o = 32'h00000000 /* 0xe0a0 */;
                14377: data_o = 32'h00000000 /* 0xe0a4 */;
                14378: data_o = 32'h00000000 /* 0xe0a8 */;
                14379: data_o = 32'h00000000 /* 0xe0ac */;
                14380: data_o = 32'h00000000 /* 0xe0b0 */;
                14381: data_o = 32'h00000000 /* 0xe0b4 */;
                14382: data_o = 32'h00000000 /* 0xe0b8 */;
                14383: data_o = 32'h00000000 /* 0xe0bc */;
                14384: data_o = 32'h00000000 /* 0xe0c0 */;
                14385: data_o = 32'h00000000 /* 0xe0c4 */;
                14386: data_o = 32'h00000000 /* 0xe0c8 */;
                14387: data_o = 32'h00000000 /* 0xe0cc */;
                14388: data_o = 32'h00000000 /* 0xe0d0 */;
                14389: data_o = 32'h00000000 /* 0xe0d4 */;
                14390: data_o = 32'h00000000 /* 0xe0d8 */;
                14391: data_o = 32'h00000000 /* 0xe0dc */;
                14392: data_o = 32'h00000000 /* 0xe0e0 */;
                14393: data_o = 32'h00000000 /* 0xe0e4 */;
                14394: data_o = 32'h00000000 /* 0xe0e8 */;
                14395: data_o = 32'h00000000 /* 0xe0ec */;
                14396: data_o = 32'h00000000 /* 0xe0f0 */;
                14397: data_o = 32'h00000000 /* 0xe0f4 */;
                14398: data_o = 32'h00000000 /* 0xe0f8 */;
                14399: data_o = 32'h00000000 /* 0xe0fc */;
                14400: data_o = 32'h00000000 /* 0xe100 */;
                14401: data_o = 32'h00000000 /* 0xe104 */;
                14402: data_o = 32'h00000000 /* 0xe108 */;
                14403: data_o = 32'h00000000 /* 0xe10c */;
                14404: data_o = 32'h00000000 /* 0xe110 */;
                14405: data_o = 32'h00000000 /* 0xe114 */;
                14406: data_o = 32'h00000000 /* 0xe118 */;
                14407: data_o = 32'h00000000 /* 0xe11c */;
                14408: data_o = 32'h00000000 /* 0xe120 */;
                14409: data_o = 32'h00000000 /* 0xe124 */;
                14410: data_o = 32'h00000000 /* 0xe128 */;
                14411: data_o = 32'h00000000 /* 0xe12c */;
                14412: data_o = 32'h00000000 /* 0xe130 */;
                14413: data_o = 32'h00000000 /* 0xe134 */;
                14414: data_o = 32'h00000000 /* 0xe138 */;
                14415: data_o = 32'h00000000 /* 0xe13c */;
                14416: data_o = 32'h00000000 /* 0xe140 */;
                14417: data_o = 32'h00000000 /* 0xe144 */;
                14418: data_o = 32'h00000000 /* 0xe148 */;
                14419: data_o = 32'h00000000 /* 0xe14c */;
                14420: data_o = 32'h00000000 /* 0xe150 */;
                14421: data_o = 32'h00000000 /* 0xe154 */;
                14422: data_o = 32'h00000000 /* 0xe158 */;
                14423: data_o = 32'h00000000 /* 0xe15c */;
                14424: data_o = 32'h00000000 /* 0xe160 */;
                14425: data_o = 32'h00000000 /* 0xe164 */;
                14426: data_o = 32'h00000000 /* 0xe168 */;
                14427: data_o = 32'h00000000 /* 0xe16c */;
                14428: data_o = 32'h00000000 /* 0xe170 */;
                14429: data_o = 32'h00000000 /* 0xe174 */;
                14430: data_o = 32'h00000000 /* 0xe178 */;
                14431: data_o = 32'h00000000 /* 0xe17c */;
                14432: data_o = 32'h00000000 /* 0xe180 */;
                14433: data_o = 32'h00000000 /* 0xe184 */;
                14434: data_o = 32'h00000000 /* 0xe188 */;
                14435: data_o = 32'h00000000 /* 0xe18c */;
                14436: data_o = 32'h00000000 /* 0xe190 */;
                14437: data_o = 32'h00000000 /* 0xe194 */;
                14438: data_o = 32'h00000000 /* 0xe198 */;
                14439: data_o = 32'h00000000 /* 0xe19c */;
                14440: data_o = 32'h00000000 /* 0xe1a0 */;
                14441: data_o = 32'h00000000 /* 0xe1a4 */;
                14442: data_o = 32'h00000000 /* 0xe1a8 */;
                14443: data_o = 32'h00000000 /* 0xe1ac */;
                14444: data_o = 32'h00000000 /* 0xe1b0 */;
                14445: data_o = 32'h00000000 /* 0xe1b4 */;
                14446: data_o = 32'h00000000 /* 0xe1b8 */;
                14447: data_o = 32'h00000000 /* 0xe1bc */;
                14448: data_o = 32'h00000000 /* 0xe1c0 */;
                14449: data_o = 32'h00000000 /* 0xe1c4 */;
                14450: data_o = 32'h00000000 /* 0xe1c8 */;
                14451: data_o = 32'h00000000 /* 0xe1cc */;
                14452: data_o = 32'h00000000 /* 0xe1d0 */;
                14453: data_o = 32'h00000000 /* 0xe1d4 */;
                14454: data_o = 32'h00000000 /* 0xe1d8 */;
                14455: data_o = 32'h00000000 /* 0xe1dc */;
                14456: data_o = 32'h00000000 /* 0xe1e0 */;
                14457: data_o = 32'h00000000 /* 0xe1e4 */;
                14458: data_o = 32'h00000000 /* 0xe1e8 */;
                14459: data_o = 32'h00000000 /* 0xe1ec */;
                14460: data_o = 32'h00000000 /* 0xe1f0 */;
                14461: data_o = 32'h00000000 /* 0xe1f4 */;
                14462: data_o = 32'h00000000 /* 0xe1f8 */;
                14463: data_o = 32'h00000000 /* 0xe1fc */;
                14464: data_o = 32'h00000000 /* 0xe200 */;
                14465: data_o = 32'h00000000 /* 0xe204 */;
                14466: data_o = 32'h00000000 /* 0xe208 */;
                14467: data_o = 32'h00000000 /* 0xe20c */;
                14468: data_o = 32'h00000000 /* 0xe210 */;
                14469: data_o = 32'h00000000 /* 0xe214 */;
                14470: data_o = 32'h00000000 /* 0xe218 */;
                14471: data_o = 32'h00000000 /* 0xe21c */;
                14472: data_o = 32'h00000000 /* 0xe220 */;
                14473: data_o = 32'h00000000 /* 0xe224 */;
                14474: data_o = 32'h00000000 /* 0xe228 */;
                14475: data_o = 32'h00000000 /* 0xe22c */;
                14476: data_o = 32'h00000000 /* 0xe230 */;
                14477: data_o = 32'h00000000 /* 0xe234 */;
                14478: data_o = 32'h00000000 /* 0xe238 */;
                14479: data_o = 32'h00000000 /* 0xe23c */;
                14480: data_o = 32'h00000000 /* 0xe240 */;
                14481: data_o = 32'h00000000 /* 0xe244 */;
                14482: data_o = 32'h00000000 /* 0xe248 */;
                14483: data_o = 32'h00000000 /* 0xe24c */;
                14484: data_o = 32'h00000000 /* 0xe250 */;
                14485: data_o = 32'h00000000 /* 0xe254 */;
                14486: data_o = 32'h00000000 /* 0xe258 */;
                14487: data_o = 32'h00000000 /* 0xe25c */;
                14488: data_o = 32'h00000000 /* 0xe260 */;
                14489: data_o = 32'h00000000 /* 0xe264 */;
                14490: data_o = 32'h00000000 /* 0xe268 */;
                14491: data_o = 32'h00000000 /* 0xe26c */;
                14492: data_o = 32'h00000000 /* 0xe270 */;
                14493: data_o = 32'h00000000 /* 0xe274 */;
                14494: data_o = 32'h00000000 /* 0xe278 */;
                14495: data_o = 32'h00000000 /* 0xe27c */;
                14496: data_o = 32'h00000000 /* 0xe280 */;
                14497: data_o = 32'h00000000 /* 0xe284 */;
                14498: data_o = 32'h00000000 /* 0xe288 */;
                14499: data_o = 32'h00000000 /* 0xe28c */;
                14500: data_o = 32'h00000000 /* 0xe290 */;
                14501: data_o = 32'h00000000 /* 0xe294 */;
                14502: data_o = 32'h00000000 /* 0xe298 */;
                14503: data_o = 32'h00000000 /* 0xe29c */;
                14504: data_o = 32'h00000000 /* 0xe2a0 */;
                14505: data_o = 32'h00000000 /* 0xe2a4 */;
                14506: data_o = 32'h00000000 /* 0xe2a8 */;
                14507: data_o = 32'h00000000 /* 0xe2ac */;
                14508: data_o = 32'h00000000 /* 0xe2b0 */;
                14509: data_o = 32'h00000000 /* 0xe2b4 */;
                14510: data_o = 32'h00000000 /* 0xe2b8 */;
                14511: data_o = 32'h00000000 /* 0xe2bc */;
                14512: data_o = 32'h00000000 /* 0xe2c0 */;
                14513: data_o = 32'h00000000 /* 0xe2c4 */;
                14514: data_o = 32'h00000000 /* 0xe2c8 */;
                14515: data_o = 32'h00000000 /* 0xe2cc */;
                14516: data_o = 32'h00000000 /* 0xe2d0 */;
                14517: data_o = 32'h00000000 /* 0xe2d4 */;
                14518: data_o = 32'h00000000 /* 0xe2d8 */;
                14519: data_o = 32'h00000000 /* 0xe2dc */;
                14520: data_o = 32'h00000000 /* 0xe2e0 */;
                14521: data_o = 32'h00000000 /* 0xe2e4 */;
                14522: data_o = 32'h00000000 /* 0xe2e8 */;
                14523: data_o = 32'h00000000 /* 0xe2ec */;
                14524: data_o = 32'h00000000 /* 0xe2f0 */;
                14525: data_o = 32'h00000000 /* 0xe2f4 */;
                14526: data_o = 32'h00000000 /* 0xe2f8 */;
                14527: data_o = 32'h00000000 /* 0xe2fc */;
                14528: data_o = 32'h00000000 /* 0xe300 */;
                14529: data_o = 32'h00000000 /* 0xe304 */;
                14530: data_o = 32'h00000000 /* 0xe308 */;
                14531: data_o = 32'h00000000 /* 0xe30c */;
                14532: data_o = 32'h00000000 /* 0xe310 */;
                14533: data_o = 32'h00000000 /* 0xe314 */;
                14534: data_o = 32'h00000000 /* 0xe318 */;
                14535: data_o = 32'h00000000 /* 0xe31c */;
                14536: data_o = 32'h00000000 /* 0xe320 */;
                14537: data_o = 32'h00000000 /* 0xe324 */;
                14538: data_o = 32'h00000000 /* 0xe328 */;
                14539: data_o = 32'h00000000 /* 0xe32c */;
                14540: data_o = 32'h00000000 /* 0xe330 */;
                14541: data_o = 32'h00000000 /* 0xe334 */;
                14542: data_o = 32'h00000000 /* 0xe338 */;
                14543: data_o = 32'h00000000 /* 0xe33c */;
                14544: data_o = 32'h00000000 /* 0xe340 */;
                14545: data_o = 32'h00000000 /* 0xe344 */;
                14546: data_o = 32'h00000000 /* 0xe348 */;
                14547: data_o = 32'h00000000 /* 0xe34c */;
                14548: data_o = 32'h00000000 /* 0xe350 */;
                14549: data_o = 32'h00000000 /* 0xe354 */;
                14550: data_o = 32'h00000000 /* 0xe358 */;
                14551: data_o = 32'h00000000 /* 0xe35c */;
                14552: data_o = 32'h00000000 /* 0xe360 */;
                14553: data_o = 32'h00000000 /* 0xe364 */;
                14554: data_o = 32'h00000000 /* 0xe368 */;
                14555: data_o = 32'h00000000 /* 0xe36c */;
                14556: data_o = 32'h00000000 /* 0xe370 */;
                14557: data_o = 32'h00000000 /* 0xe374 */;
                14558: data_o = 32'h00000000 /* 0xe378 */;
                14559: data_o = 32'h00000000 /* 0xe37c */;
                14560: data_o = 32'h00000000 /* 0xe380 */;
                14561: data_o = 32'h00000000 /* 0xe384 */;
                14562: data_o = 32'h00000000 /* 0xe388 */;
                14563: data_o = 32'h00000000 /* 0xe38c */;
                14564: data_o = 32'h00000000 /* 0xe390 */;
                14565: data_o = 32'h00000000 /* 0xe394 */;
                14566: data_o = 32'h00000000 /* 0xe398 */;
                14567: data_o = 32'h00000000 /* 0xe39c */;
                14568: data_o = 32'h00000000 /* 0xe3a0 */;
                14569: data_o = 32'h00000000 /* 0xe3a4 */;
                14570: data_o = 32'h00000000 /* 0xe3a8 */;
                14571: data_o = 32'h00000000 /* 0xe3ac */;
                14572: data_o = 32'h00000000 /* 0xe3b0 */;
                14573: data_o = 32'h00000000 /* 0xe3b4 */;
                14574: data_o = 32'h00000000 /* 0xe3b8 */;
                14575: data_o = 32'h00000000 /* 0xe3bc */;
                14576: data_o = 32'h00000000 /* 0xe3c0 */;
                14577: data_o = 32'h00000000 /* 0xe3c4 */;
                14578: data_o = 32'h00000000 /* 0xe3c8 */;
                14579: data_o = 32'h00000000 /* 0xe3cc */;
                14580: data_o = 32'h00000000 /* 0xe3d0 */;
                14581: data_o = 32'h00000000 /* 0xe3d4 */;
                14582: data_o = 32'h00000000 /* 0xe3d8 */;
                14583: data_o = 32'h00000000 /* 0xe3dc */;
                14584: data_o = 32'h00000000 /* 0xe3e0 */;
                14585: data_o = 32'h00000000 /* 0xe3e4 */;
                14586: data_o = 32'h00000000 /* 0xe3e8 */;
                14587: data_o = 32'h00000000 /* 0xe3ec */;
                14588: data_o = 32'h00000000 /* 0xe3f0 */;
                14589: data_o = 32'h00000000 /* 0xe3f4 */;
                14590: data_o = 32'h00000000 /* 0xe3f8 */;
                14591: data_o = 32'h00000000 /* 0xe3fc */;
                14592: data_o = 32'h00000000 /* 0xe400 */;
                14593: data_o = 32'h00000000 /* 0xe404 */;
                14594: data_o = 32'h00000000 /* 0xe408 */;
                14595: data_o = 32'h00000000 /* 0xe40c */;
                14596: data_o = 32'h00000000 /* 0xe410 */;
                14597: data_o = 32'h00000000 /* 0xe414 */;
                14598: data_o = 32'h00000000 /* 0xe418 */;
                14599: data_o = 32'h00000000 /* 0xe41c */;
                14600: data_o = 32'h00000000 /* 0xe420 */;
                14601: data_o = 32'h00000000 /* 0xe424 */;
                14602: data_o = 32'h00000000 /* 0xe428 */;
                14603: data_o = 32'h00000000 /* 0xe42c */;
                14604: data_o = 32'h00000000 /* 0xe430 */;
                14605: data_o = 32'h00000000 /* 0xe434 */;
                14606: data_o = 32'h00000000 /* 0xe438 */;
                14607: data_o = 32'h00000000 /* 0xe43c */;
                14608: data_o = 32'h00000000 /* 0xe440 */;
                14609: data_o = 32'h00000000 /* 0xe444 */;
                14610: data_o = 32'h00000000 /* 0xe448 */;
                14611: data_o = 32'h00000000 /* 0xe44c */;
                14612: data_o = 32'h00000000 /* 0xe450 */;
                14613: data_o = 32'h00000000 /* 0xe454 */;
                14614: data_o = 32'h00000000 /* 0xe458 */;
                14615: data_o = 32'h00000000 /* 0xe45c */;
                14616: data_o = 32'h00000000 /* 0xe460 */;
                14617: data_o = 32'h00000000 /* 0xe464 */;
                14618: data_o = 32'h00000000 /* 0xe468 */;
                14619: data_o = 32'h00000000 /* 0xe46c */;
                14620: data_o = 32'h00000000 /* 0xe470 */;
                14621: data_o = 32'h00000000 /* 0xe474 */;
                14622: data_o = 32'h00000000 /* 0xe478 */;
                14623: data_o = 32'h00000000 /* 0xe47c */;
                14624: data_o = 32'h00000000 /* 0xe480 */;
                14625: data_o = 32'h00000000 /* 0xe484 */;
                14626: data_o = 32'h00000000 /* 0xe488 */;
                14627: data_o = 32'h00000000 /* 0xe48c */;
                14628: data_o = 32'h00000000 /* 0xe490 */;
                14629: data_o = 32'h00000000 /* 0xe494 */;
                14630: data_o = 32'h00000000 /* 0xe498 */;
                14631: data_o = 32'h00000000 /* 0xe49c */;
                14632: data_o = 32'h00000000 /* 0xe4a0 */;
                14633: data_o = 32'h00000000 /* 0xe4a4 */;
                14634: data_o = 32'h00000000 /* 0xe4a8 */;
                14635: data_o = 32'h00000000 /* 0xe4ac */;
                14636: data_o = 32'h00000000 /* 0xe4b0 */;
                14637: data_o = 32'h00000000 /* 0xe4b4 */;
                14638: data_o = 32'h00000000 /* 0xe4b8 */;
                14639: data_o = 32'h00000000 /* 0xe4bc */;
                14640: data_o = 32'h00000000 /* 0xe4c0 */;
                14641: data_o = 32'h00000000 /* 0xe4c4 */;
                14642: data_o = 32'h00000000 /* 0xe4c8 */;
                14643: data_o = 32'h00000000 /* 0xe4cc */;
                14644: data_o = 32'h00000000 /* 0xe4d0 */;
                14645: data_o = 32'h00000000 /* 0xe4d4 */;
                14646: data_o = 32'h00000000 /* 0xe4d8 */;
                14647: data_o = 32'h00000000 /* 0xe4dc */;
                14648: data_o = 32'h00000000 /* 0xe4e0 */;
                14649: data_o = 32'h00000000 /* 0xe4e4 */;
                14650: data_o = 32'h00000000 /* 0xe4e8 */;
                14651: data_o = 32'h00000000 /* 0xe4ec */;
                14652: data_o = 32'h00000000 /* 0xe4f0 */;
                14653: data_o = 32'h00000000 /* 0xe4f4 */;
                14654: data_o = 32'h00000000 /* 0xe4f8 */;
                14655: data_o = 32'h00000000 /* 0xe4fc */;
                14656: data_o = 32'h00000000 /* 0xe500 */;
                14657: data_o = 32'h00000000 /* 0xe504 */;
                14658: data_o = 32'h00000000 /* 0xe508 */;
                14659: data_o = 32'h00000000 /* 0xe50c */;
                14660: data_o = 32'h00000000 /* 0xe510 */;
                14661: data_o = 32'h00000000 /* 0xe514 */;
                14662: data_o = 32'h00000000 /* 0xe518 */;
                14663: data_o = 32'h00000000 /* 0xe51c */;
                14664: data_o = 32'h00000000 /* 0xe520 */;
                14665: data_o = 32'h00000000 /* 0xe524 */;
                14666: data_o = 32'h00000000 /* 0xe528 */;
                14667: data_o = 32'h00000000 /* 0xe52c */;
                14668: data_o = 32'h00000000 /* 0xe530 */;
                14669: data_o = 32'h00000000 /* 0xe534 */;
                14670: data_o = 32'h00000000 /* 0xe538 */;
                14671: data_o = 32'h00000000 /* 0xe53c */;
                14672: data_o = 32'h00000000 /* 0xe540 */;
                14673: data_o = 32'h00000000 /* 0xe544 */;
                14674: data_o = 32'h00000000 /* 0xe548 */;
                14675: data_o = 32'h00000000 /* 0xe54c */;
                14676: data_o = 32'h00000000 /* 0xe550 */;
                14677: data_o = 32'h00000000 /* 0xe554 */;
                14678: data_o = 32'h00000000 /* 0xe558 */;
                14679: data_o = 32'h00000000 /* 0xe55c */;
                14680: data_o = 32'h00000000 /* 0xe560 */;
                14681: data_o = 32'h00000000 /* 0xe564 */;
                14682: data_o = 32'h00000000 /* 0xe568 */;
                14683: data_o = 32'h00000000 /* 0xe56c */;
                14684: data_o = 32'h00000000 /* 0xe570 */;
                14685: data_o = 32'h00000000 /* 0xe574 */;
                14686: data_o = 32'h00000000 /* 0xe578 */;
                14687: data_o = 32'h00000000 /* 0xe57c */;
                14688: data_o = 32'h00000000 /* 0xe580 */;
                14689: data_o = 32'h00000000 /* 0xe584 */;
                14690: data_o = 32'h00000000 /* 0xe588 */;
                14691: data_o = 32'h00000000 /* 0xe58c */;
                14692: data_o = 32'h00000000 /* 0xe590 */;
                14693: data_o = 32'h00000000 /* 0xe594 */;
                14694: data_o = 32'h00000000 /* 0xe598 */;
                14695: data_o = 32'h00000000 /* 0xe59c */;
                14696: data_o = 32'h00000000 /* 0xe5a0 */;
                14697: data_o = 32'h00000000 /* 0xe5a4 */;
                14698: data_o = 32'h00000000 /* 0xe5a8 */;
                14699: data_o = 32'h00000000 /* 0xe5ac */;
                14700: data_o = 32'h00000000 /* 0xe5b0 */;
                14701: data_o = 32'h00000000 /* 0xe5b4 */;
                14702: data_o = 32'h00000000 /* 0xe5b8 */;
                14703: data_o = 32'h00000000 /* 0xe5bc */;
                14704: data_o = 32'h00000000 /* 0xe5c0 */;
                14705: data_o = 32'h00000000 /* 0xe5c4 */;
                14706: data_o = 32'h00000000 /* 0xe5c8 */;
                14707: data_o = 32'h00000000 /* 0xe5cc */;
                14708: data_o = 32'h00000000 /* 0xe5d0 */;
                14709: data_o = 32'h00000000 /* 0xe5d4 */;
                14710: data_o = 32'h00000000 /* 0xe5d8 */;
                14711: data_o = 32'h00000000 /* 0xe5dc */;
                14712: data_o = 32'h00000000 /* 0xe5e0 */;
                14713: data_o = 32'h00000000 /* 0xe5e4 */;
                14714: data_o = 32'h00000000 /* 0xe5e8 */;
                14715: data_o = 32'h00000000 /* 0xe5ec */;
                14716: data_o = 32'h00000000 /* 0xe5f0 */;
                14717: data_o = 32'h00000000 /* 0xe5f4 */;
                14718: data_o = 32'h00000000 /* 0xe5f8 */;
                14719: data_o = 32'h00000000 /* 0xe5fc */;
                14720: data_o = 32'h00000000 /* 0xe600 */;
                14721: data_o = 32'h00000000 /* 0xe604 */;
                14722: data_o = 32'h00000000 /* 0xe608 */;
                14723: data_o = 32'h00000000 /* 0xe60c */;
                14724: data_o = 32'h00000000 /* 0xe610 */;
                14725: data_o = 32'h00000000 /* 0xe614 */;
                14726: data_o = 32'h00000000 /* 0xe618 */;
                14727: data_o = 32'h00000000 /* 0xe61c */;
                14728: data_o = 32'h00000000 /* 0xe620 */;
                14729: data_o = 32'h00000000 /* 0xe624 */;
                14730: data_o = 32'h00000000 /* 0xe628 */;
                14731: data_o = 32'h00000000 /* 0xe62c */;
                14732: data_o = 32'h00000000 /* 0xe630 */;
                14733: data_o = 32'h00000000 /* 0xe634 */;
                14734: data_o = 32'h00000000 /* 0xe638 */;
                14735: data_o = 32'h00000000 /* 0xe63c */;
                14736: data_o = 32'h00000000 /* 0xe640 */;
                14737: data_o = 32'h00000000 /* 0xe644 */;
                14738: data_o = 32'h00000000 /* 0xe648 */;
                14739: data_o = 32'h00000000 /* 0xe64c */;
                14740: data_o = 32'h00000000 /* 0xe650 */;
                14741: data_o = 32'h00000000 /* 0xe654 */;
                14742: data_o = 32'h00000000 /* 0xe658 */;
                14743: data_o = 32'h00000000 /* 0xe65c */;
                14744: data_o = 32'h00000000 /* 0xe660 */;
                14745: data_o = 32'h00000000 /* 0xe664 */;
                14746: data_o = 32'h00000000 /* 0xe668 */;
                14747: data_o = 32'h00000000 /* 0xe66c */;
                14748: data_o = 32'h00000000 /* 0xe670 */;
                14749: data_o = 32'h00000000 /* 0xe674 */;
                14750: data_o = 32'h00000000 /* 0xe678 */;
                14751: data_o = 32'h00000000 /* 0xe67c */;
                14752: data_o = 32'h00000000 /* 0xe680 */;
                14753: data_o = 32'h00000000 /* 0xe684 */;
                14754: data_o = 32'h00000000 /* 0xe688 */;
                14755: data_o = 32'h00000000 /* 0xe68c */;
                14756: data_o = 32'h00000000 /* 0xe690 */;
                14757: data_o = 32'h00000000 /* 0xe694 */;
                14758: data_o = 32'h00000000 /* 0xe698 */;
                14759: data_o = 32'h00000000 /* 0xe69c */;
                14760: data_o = 32'h00000000 /* 0xe6a0 */;
                14761: data_o = 32'h00000000 /* 0xe6a4 */;
                14762: data_o = 32'h00000000 /* 0xe6a8 */;
                14763: data_o = 32'h00000000 /* 0xe6ac */;
                14764: data_o = 32'h00000000 /* 0xe6b0 */;
                14765: data_o = 32'h00000000 /* 0xe6b4 */;
                14766: data_o = 32'h00000000 /* 0xe6b8 */;
                14767: data_o = 32'h00000000 /* 0xe6bc */;
                14768: data_o = 32'h00000000 /* 0xe6c0 */;
                14769: data_o = 32'h00000000 /* 0xe6c4 */;
                14770: data_o = 32'h00000000 /* 0xe6c8 */;
                14771: data_o = 32'h00000000 /* 0xe6cc */;
                14772: data_o = 32'h00000000 /* 0xe6d0 */;
                14773: data_o = 32'h00000000 /* 0xe6d4 */;
                14774: data_o = 32'h00000000 /* 0xe6d8 */;
                14775: data_o = 32'h00000000 /* 0xe6dc */;
                14776: data_o = 32'h00000000 /* 0xe6e0 */;
                14777: data_o = 32'h00000000 /* 0xe6e4 */;
                14778: data_o = 32'h00000000 /* 0xe6e8 */;
                14779: data_o = 32'h00000000 /* 0xe6ec */;
                14780: data_o = 32'h00000000 /* 0xe6f0 */;
                14781: data_o = 32'h00000000 /* 0xe6f4 */;
                14782: data_o = 32'h00000000 /* 0xe6f8 */;
                14783: data_o = 32'h00000000 /* 0xe6fc */;
                14784: data_o = 32'h00000000 /* 0xe700 */;
                14785: data_o = 32'h00000000 /* 0xe704 */;
                14786: data_o = 32'h00000000 /* 0xe708 */;
                14787: data_o = 32'h00000000 /* 0xe70c */;
                14788: data_o = 32'h00000000 /* 0xe710 */;
                14789: data_o = 32'h00000000 /* 0xe714 */;
                14790: data_o = 32'h00000000 /* 0xe718 */;
                14791: data_o = 32'h00000000 /* 0xe71c */;
                14792: data_o = 32'h00000000 /* 0xe720 */;
                14793: data_o = 32'h00000000 /* 0xe724 */;
                14794: data_o = 32'h00000000 /* 0xe728 */;
                14795: data_o = 32'h00000000 /* 0xe72c */;
                14796: data_o = 32'h00000000 /* 0xe730 */;
                14797: data_o = 32'h00000000 /* 0xe734 */;
                14798: data_o = 32'h00000000 /* 0xe738 */;
                14799: data_o = 32'h00000000 /* 0xe73c */;
                14800: data_o = 32'h00000000 /* 0xe740 */;
                14801: data_o = 32'h00000000 /* 0xe744 */;
                14802: data_o = 32'h00000000 /* 0xe748 */;
                14803: data_o = 32'h00000000 /* 0xe74c */;
                14804: data_o = 32'h00000000 /* 0xe750 */;
                14805: data_o = 32'h00000000 /* 0xe754 */;
                14806: data_o = 32'h00000000 /* 0xe758 */;
                14807: data_o = 32'h00000000 /* 0xe75c */;
                14808: data_o = 32'h00000000 /* 0xe760 */;
                14809: data_o = 32'h00000000 /* 0xe764 */;
                14810: data_o = 32'h00000000 /* 0xe768 */;
                14811: data_o = 32'h00000000 /* 0xe76c */;
                14812: data_o = 32'h00000000 /* 0xe770 */;
                14813: data_o = 32'h00000000 /* 0xe774 */;
                14814: data_o = 32'h00000000 /* 0xe778 */;
                14815: data_o = 32'h00000000 /* 0xe77c */;
                14816: data_o = 32'h00000000 /* 0xe780 */;
                14817: data_o = 32'h00000000 /* 0xe784 */;
                14818: data_o = 32'h00000000 /* 0xe788 */;
                14819: data_o = 32'h00000000 /* 0xe78c */;
                14820: data_o = 32'h00000000 /* 0xe790 */;
                14821: data_o = 32'h00000000 /* 0xe794 */;
                14822: data_o = 32'h00000000 /* 0xe798 */;
                14823: data_o = 32'h00000000 /* 0xe79c */;
                14824: data_o = 32'h00000000 /* 0xe7a0 */;
                14825: data_o = 32'h00000000 /* 0xe7a4 */;
                14826: data_o = 32'h00000000 /* 0xe7a8 */;
                14827: data_o = 32'h00000000 /* 0xe7ac */;
                14828: data_o = 32'h00000000 /* 0xe7b0 */;
                14829: data_o = 32'h00000000 /* 0xe7b4 */;
                14830: data_o = 32'h00000000 /* 0xe7b8 */;
                14831: data_o = 32'h00000000 /* 0xe7bc */;
                14832: data_o = 32'h00000000 /* 0xe7c0 */;
                14833: data_o = 32'h00000000 /* 0xe7c4 */;
                14834: data_o = 32'h00000000 /* 0xe7c8 */;
                14835: data_o = 32'h00000000 /* 0xe7cc */;
                14836: data_o = 32'h00000000 /* 0xe7d0 */;
                14837: data_o = 32'h00000000 /* 0xe7d4 */;
                14838: data_o = 32'h00000000 /* 0xe7d8 */;
                14839: data_o = 32'h00000000 /* 0xe7dc */;
                14840: data_o = 32'h00000000 /* 0xe7e0 */;
                14841: data_o = 32'h00000000 /* 0xe7e4 */;
                14842: data_o = 32'h00000000 /* 0xe7e8 */;
                14843: data_o = 32'h00000000 /* 0xe7ec */;
                14844: data_o = 32'h00000000 /* 0xe7f0 */;
                14845: data_o = 32'h00000000 /* 0xe7f4 */;
                14846: data_o = 32'h00000000 /* 0xe7f8 */;
                14847: data_o = 32'h00000000 /* 0xe7fc */;
                14848: data_o = 32'h00000000 /* 0xe800 */;
                14849: data_o = 32'h00000000 /* 0xe804 */;
                14850: data_o = 32'h00000000 /* 0xe808 */;
                14851: data_o = 32'h00000000 /* 0xe80c */;
                14852: data_o = 32'h00000000 /* 0xe810 */;
                14853: data_o = 32'h00000000 /* 0xe814 */;
                14854: data_o = 32'h00000000 /* 0xe818 */;
                14855: data_o = 32'h00000000 /* 0xe81c */;
                14856: data_o = 32'h00000000 /* 0xe820 */;
                14857: data_o = 32'h00000000 /* 0xe824 */;
                14858: data_o = 32'h00000000 /* 0xe828 */;
                14859: data_o = 32'h00000000 /* 0xe82c */;
                14860: data_o = 32'h00000000 /* 0xe830 */;
                14861: data_o = 32'h00000000 /* 0xe834 */;
                14862: data_o = 32'h00000000 /* 0xe838 */;
                14863: data_o = 32'h00000000 /* 0xe83c */;
                14864: data_o = 32'h00000000 /* 0xe840 */;
                14865: data_o = 32'h00000000 /* 0xe844 */;
                14866: data_o = 32'h00000000 /* 0xe848 */;
                14867: data_o = 32'h00000000 /* 0xe84c */;
                14868: data_o = 32'h00000000 /* 0xe850 */;
                14869: data_o = 32'h00000000 /* 0xe854 */;
                14870: data_o = 32'h00000000 /* 0xe858 */;
                14871: data_o = 32'h00000000 /* 0xe85c */;
                14872: data_o = 32'h00000000 /* 0xe860 */;
                14873: data_o = 32'h00000000 /* 0xe864 */;
                14874: data_o = 32'h00000000 /* 0xe868 */;
                14875: data_o = 32'h00000000 /* 0xe86c */;
                14876: data_o = 32'h00000000 /* 0xe870 */;
                14877: data_o = 32'h00000000 /* 0xe874 */;
                14878: data_o = 32'h00000000 /* 0xe878 */;
                14879: data_o = 32'h00000000 /* 0xe87c */;
                14880: data_o = 32'h00000000 /* 0xe880 */;
                14881: data_o = 32'h00000000 /* 0xe884 */;
                14882: data_o = 32'h00000000 /* 0xe888 */;
                14883: data_o = 32'h00000000 /* 0xe88c */;
                14884: data_o = 32'h00000000 /* 0xe890 */;
                14885: data_o = 32'h00000000 /* 0xe894 */;
                14886: data_o = 32'h00000000 /* 0xe898 */;
                14887: data_o = 32'h00000000 /* 0xe89c */;
                14888: data_o = 32'h00000000 /* 0xe8a0 */;
                14889: data_o = 32'h00000000 /* 0xe8a4 */;
                14890: data_o = 32'h00000000 /* 0xe8a8 */;
                14891: data_o = 32'h00000000 /* 0xe8ac */;
                14892: data_o = 32'h00000000 /* 0xe8b0 */;
                14893: data_o = 32'h00000000 /* 0xe8b4 */;
                14894: data_o = 32'h00000000 /* 0xe8b8 */;
                14895: data_o = 32'h00000000 /* 0xe8bc */;
                14896: data_o = 32'h00000000 /* 0xe8c0 */;
                14897: data_o = 32'h00000000 /* 0xe8c4 */;
                14898: data_o = 32'h00000000 /* 0xe8c8 */;
                14899: data_o = 32'h00000000 /* 0xe8cc */;
                14900: data_o = 32'h00000000 /* 0xe8d0 */;
                14901: data_o = 32'h00000000 /* 0xe8d4 */;
                14902: data_o = 32'h00000000 /* 0xe8d8 */;
                14903: data_o = 32'h00000000 /* 0xe8dc */;
                14904: data_o = 32'h00000000 /* 0xe8e0 */;
                14905: data_o = 32'h00000000 /* 0xe8e4 */;
                14906: data_o = 32'h00000000 /* 0xe8e8 */;
                14907: data_o = 32'h00000000 /* 0xe8ec */;
                14908: data_o = 32'h00000000 /* 0xe8f0 */;
                14909: data_o = 32'h00000000 /* 0xe8f4 */;
                14910: data_o = 32'h00000000 /* 0xe8f8 */;
                14911: data_o = 32'h00000000 /* 0xe8fc */;
                14912: data_o = 32'h00000000 /* 0xe900 */;
                14913: data_o = 32'h00000000 /* 0xe904 */;
                14914: data_o = 32'h00000000 /* 0xe908 */;
                14915: data_o = 32'h00000000 /* 0xe90c */;
                14916: data_o = 32'h00000000 /* 0xe910 */;
                14917: data_o = 32'h00000000 /* 0xe914 */;
                14918: data_o = 32'h00000000 /* 0xe918 */;
                14919: data_o = 32'h00000000 /* 0xe91c */;
                14920: data_o = 32'h00000000 /* 0xe920 */;
                14921: data_o = 32'h00000000 /* 0xe924 */;
                14922: data_o = 32'h00000000 /* 0xe928 */;
                14923: data_o = 32'h00000000 /* 0xe92c */;
                14924: data_o = 32'h00000000 /* 0xe930 */;
                14925: data_o = 32'h00000000 /* 0xe934 */;
                14926: data_o = 32'h00000000 /* 0xe938 */;
                14927: data_o = 32'h00000000 /* 0xe93c */;
                14928: data_o = 32'h00000000 /* 0xe940 */;
                14929: data_o = 32'h00000000 /* 0xe944 */;
                14930: data_o = 32'h00000000 /* 0xe948 */;
                14931: data_o = 32'h00000000 /* 0xe94c */;
                14932: data_o = 32'h00000000 /* 0xe950 */;
                14933: data_o = 32'h00000000 /* 0xe954 */;
                14934: data_o = 32'h00000000 /* 0xe958 */;
                14935: data_o = 32'h00000000 /* 0xe95c */;
                14936: data_o = 32'h00000000 /* 0xe960 */;
                14937: data_o = 32'h00000000 /* 0xe964 */;
                14938: data_o = 32'h00000000 /* 0xe968 */;
                14939: data_o = 32'h00000000 /* 0xe96c */;
                14940: data_o = 32'h00000000 /* 0xe970 */;
                14941: data_o = 32'h00000000 /* 0xe974 */;
                14942: data_o = 32'h00000000 /* 0xe978 */;
                14943: data_o = 32'h00000000 /* 0xe97c */;
                14944: data_o = 32'h00000000 /* 0xe980 */;
                14945: data_o = 32'h00000000 /* 0xe984 */;
                14946: data_o = 32'h00000000 /* 0xe988 */;
                14947: data_o = 32'h00000000 /* 0xe98c */;
                14948: data_o = 32'h00000000 /* 0xe990 */;
                14949: data_o = 32'h00000000 /* 0xe994 */;
                14950: data_o = 32'h00000000 /* 0xe998 */;
                14951: data_o = 32'h00000000 /* 0xe99c */;
                14952: data_o = 32'h00000000 /* 0xe9a0 */;
                14953: data_o = 32'h00000000 /* 0xe9a4 */;
                14954: data_o = 32'h00000000 /* 0xe9a8 */;
                14955: data_o = 32'h00000000 /* 0xe9ac */;
                14956: data_o = 32'h00000000 /* 0xe9b0 */;
                14957: data_o = 32'h00000000 /* 0xe9b4 */;
                14958: data_o = 32'h00000000 /* 0xe9b8 */;
                14959: data_o = 32'h00000000 /* 0xe9bc */;
                14960: data_o = 32'h00000000 /* 0xe9c0 */;
                14961: data_o = 32'h00000000 /* 0xe9c4 */;
                14962: data_o = 32'h00000000 /* 0xe9c8 */;
                14963: data_o = 32'h00000000 /* 0xe9cc */;
                14964: data_o = 32'h00000000 /* 0xe9d0 */;
                14965: data_o = 32'h00000000 /* 0xe9d4 */;
                14966: data_o = 32'h00000000 /* 0xe9d8 */;
                14967: data_o = 32'h00000000 /* 0xe9dc */;
                14968: data_o = 32'h00000000 /* 0xe9e0 */;
                14969: data_o = 32'h00000000 /* 0xe9e4 */;
                14970: data_o = 32'h00000000 /* 0xe9e8 */;
                14971: data_o = 32'h00000000 /* 0xe9ec */;
                14972: data_o = 32'h00000000 /* 0xe9f0 */;
                14973: data_o = 32'h00000000 /* 0xe9f4 */;
                14974: data_o = 32'h00000000 /* 0xe9f8 */;
                14975: data_o = 32'h00000000 /* 0xe9fc */;
                14976: data_o = 32'h00000000 /* 0xea00 */;
                14977: data_o = 32'h00000000 /* 0xea04 */;
                14978: data_o = 32'h00000000 /* 0xea08 */;
                14979: data_o = 32'h00000000 /* 0xea0c */;
                14980: data_o = 32'h00000000 /* 0xea10 */;
                14981: data_o = 32'h00000000 /* 0xea14 */;
                14982: data_o = 32'h00000000 /* 0xea18 */;
                14983: data_o = 32'h00000000 /* 0xea1c */;
                14984: data_o = 32'h00000000 /* 0xea20 */;
                14985: data_o = 32'h00000000 /* 0xea24 */;
                14986: data_o = 32'h00000000 /* 0xea28 */;
                14987: data_o = 32'h00000000 /* 0xea2c */;
                14988: data_o = 32'h00000000 /* 0xea30 */;
                14989: data_o = 32'h00000000 /* 0xea34 */;
                14990: data_o = 32'h00000000 /* 0xea38 */;
                14991: data_o = 32'h00000000 /* 0xea3c */;
                14992: data_o = 32'h00000000 /* 0xea40 */;
                14993: data_o = 32'h00000000 /* 0xea44 */;
                14994: data_o = 32'h00000000 /* 0xea48 */;
                14995: data_o = 32'h00000000 /* 0xea4c */;
                14996: data_o = 32'h00000000 /* 0xea50 */;
                14997: data_o = 32'h00000000 /* 0xea54 */;
                14998: data_o = 32'h00000000 /* 0xea58 */;
                14999: data_o = 32'h00000000 /* 0xea5c */;
                15000: data_o = 32'h00000000 /* 0xea60 */;
                15001: data_o = 32'h00000000 /* 0xea64 */;
                15002: data_o = 32'h00000000 /* 0xea68 */;
                15003: data_o = 32'h00000000 /* 0xea6c */;
                15004: data_o = 32'h00000000 /* 0xea70 */;
                15005: data_o = 32'h00000000 /* 0xea74 */;
                15006: data_o = 32'h00000000 /* 0xea78 */;
                15007: data_o = 32'h00000000 /* 0xea7c */;
                15008: data_o = 32'h00000000 /* 0xea80 */;
                15009: data_o = 32'h00000000 /* 0xea84 */;
                15010: data_o = 32'h00000000 /* 0xea88 */;
                15011: data_o = 32'h00000000 /* 0xea8c */;
                15012: data_o = 32'h00000000 /* 0xea90 */;
                15013: data_o = 32'h00000000 /* 0xea94 */;
                15014: data_o = 32'h00000000 /* 0xea98 */;
                15015: data_o = 32'h00000000 /* 0xea9c */;
                15016: data_o = 32'h00000000 /* 0xeaa0 */;
                15017: data_o = 32'h00000000 /* 0xeaa4 */;
                15018: data_o = 32'h00000000 /* 0xeaa8 */;
                15019: data_o = 32'h00000000 /* 0xeaac */;
                15020: data_o = 32'h00000000 /* 0xeab0 */;
                15021: data_o = 32'h00000000 /* 0xeab4 */;
                15022: data_o = 32'h00000000 /* 0xeab8 */;
                15023: data_o = 32'h00000000 /* 0xeabc */;
                15024: data_o = 32'h00000000 /* 0xeac0 */;
                15025: data_o = 32'h00000000 /* 0xeac4 */;
                15026: data_o = 32'h00000000 /* 0xeac8 */;
                15027: data_o = 32'h00000000 /* 0xeacc */;
                15028: data_o = 32'h00000000 /* 0xead0 */;
                15029: data_o = 32'h00000000 /* 0xead4 */;
                15030: data_o = 32'h00000000 /* 0xead8 */;
                15031: data_o = 32'h00000000 /* 0xeadc */;
                15032: data_o = 32'h00000000 /* 0xeae0 */;
                15033: data_o = 32'h00000000 /* 0xeae4 */;
                15034: data_o = 32'h00000000 /* 0xeae8 */;
                15035: data_o = 32'h00000000 /* 0xeaec */;
                15036: data_o = 32'h00000000 /* 0xeaf0 */;
                15037: data_o = 32'h00000000 /* 0xeaf4 */;
                15038: data_o = 32'h00000000 /* 0xeaf8 */;
                15039: data_o = 32'h00000000 /* 0xeafc */;
                15040: data_o = 32'h00000000 /* 0xeb00 */;
                15041: data_o = 32'h00000000 /* 0xeb04 */;
                15042: data_o = 32'h00000000 /* 0xeb08 */;
                15043: data_o = 32'h00000000 /* 0xeb0c */;
                15044: data_o = 32'h00000000 /* 0xeb10 */;
                15045: data_o = 32'h00000000 /* 0xeb14 */;
                15046: data_o = 32'h00000000 /* 0xeb18 */;
                15047: data_o = 32'h00000000 /* 0xeb1c */;
                15048: data_o = 32'h00000000 /* 0xeb20 */;
                15049: data_o = 32'h00000000 /* 0xeb24 */;
                15050: data_o = 32'h00000000 /* 0xeb28 */;
                15051: data_o = 32'h00000000 /* 0xeb2c */;
                15052: data_o = 32'h00000000 /* 0xeb30 */;
                15053: data_o = 32'h00000000 /* 0xeb34 */;
                15054: data_o = 32'h00000000 /* 0xeb38 */;
                15055: data_o = 32'h00000000 /* 0xeb3c */;
                15056: data_o = 32'h00000000 /* 0xeb40 */;
                15057: data_o = 32'h00000000 /* 0xeb44 */;
                15058: data_o = 32'h00000000 /* 0xeb48 */;
                15059: data_o = 32'h00000000 /* 0xeb4c */;
                15060: data_o = 32'h00000000 /* 0xeb50 */;
                15061: data_o = 32'h00000000 /* 0xeb54 */;
                15062: data_o = 32'h00000000 /* 0xeb58 */;
                15063: data_o = 32'h00000000 /* 0xeb5c */;
                15064: data_o = 32'h00000000 /* 0xeb60 */;
                15065: data_o = 32'h00000000 /* 0xeb64 */;
                15066: data_o = 32'h00000000 /* 0xeb68 */;
                15067: data_o = 32'h00000000 /* 0xeb6c */;
                15068: data_o = 32'h00000000 /* 0xeb70 */;
                15069: data_o = 32'h00000000 /* 0xeb74 */;
                15070: data_o = 32'h00000000 /* 0xeb78 */;
                15071: data_o = 32'h00000000 /* 0xeb7c */;
                15072: data_o = 32'h00000000 /* 0xeb80 */;
                15073: data_o = 32'h00000000 /* 0xeb84 */;
                15074: data_o = 32'h00000000 /* 0xeb88 */;
                15075: data_o = 32'h00000000 /* 0xeb8c */;
                15076: data_o = 32'h00000000 /* 0xeb90 */;
                15077: data_o = 32'h00000000 /* 0xeb94 */;
                15078: data_o = 32'h00000000 /* 0xeb98 */;
                15079: data_o = 32'h00000000 /* 0xeb9c */;
                15080: data_o = 32'h00000000 /* 0xeba0 */;
                15081: data_o = 32'h00000000 /* 0xeba4 */;
                15082: data_o = 32'h00000000 /* 0xeba8 */;
                15083: data_o = 32'h00000000 /* 0xebac */;
                15084: data_o = 32'h00000000 /* 0xebb0 */;
                15085: data_o = 32'h00000000 /* 0xebb4 */;
                15086: data_o = 32'h00000000 /* 0xebb8 */;
                15087: data_o = 32'h00000000 /* 0xebbc */;
                15088: data_o = 32'h00000000 /* 0xebc0 */;
                15089: data_o = 32'h00000000 /* 0xebc4 */;
                15090: data_o = 32'h00000000 /* 0xebc8 */;
                15091: data_o = 32'h00000000 /* 0xebcc */;
                15092: data_o = 32'h00000000 /* 0xebd0 */;
                15093: data_o = 32'h00000000 /* 0xebd4 */;
                15094: data_o = 32'h00000000 /* 0xebd8 */;
                15095: data_o = 32'h00000000 /* 0xebdc */;
                15096: data_o = 32'h00000000 /* 0xebe0 */;
                15097: data_o = 32'h00000000 /* 0xebe4 */;
                15098: data_o = 32'h00000000 /* 0xebe8 */;
                15099: data_o = 32'h00000000 /* 0xebec */;
                15100: data_o = 32'h00000000 /* 0xebf0 */;
                15101: data_o = 32'h00000000 /* 0xebf4 */;
                15102: data_o = 32'h00000000 /* 0xebf8 */;
                15103: data_o = 32'h00000000 /* 0xebfc */;
                15104: data_o = 32'h00000000 /* 0xec00 */;
                15105: data_o = 32'h00000000 /* 0xec04 */;
                15106: data_o = 32'h00000000 /* 0xec08 */;
                15107: data_o = 32'h00000000 /* 0xec0c */;
                15108: data_o = 32'h00000000 /* 0xec10 */;
                15109: data_o = 32'h00000000 /* 0xec14 */;
                15110: data_o = 32'h00000000 /* 0xec18 */;
                15111: data_o = 32'h00000000 /* 0xec1c */;
                15112: data_o = 32'h00000000 /* 0xec20 */;
                15113: data_o = 32'h00000000 /* 0xec24 */;
                15114: data_o = 32'h00000000 /* 0xec28 */;
                15115: data_o = 32'h00000000 /* 0xec2c */;
                15116: data_o = 32'h00000000 /* 0xec30 */;
                15117: data_o = 32'h00000000 /* 0xec34 */;
                15118: data_o = 32'h00000000 /* 0xec38 */;
                15119: data_o = 32'h00000000 /* 0xec3c */;
                15120: data_o = 32'h00000000 /* 0xec40 */;
                15121: data_o = 32'h00000000 /* 0xec44 */;
                15122: data_o = 32'h00000000 /* 0xec48 */;
                15123: data_o = 32'h00000000 /* 0xec4c */;
                15124: data_o = 32'h00000000 /* 0xec50 */;
                15125: data_o = 32'h00000000 /* 0xec54 */;
                15126: data_o = 32'h00000000 /* 0xec58 */;
                15127: data_o = 32'h00000000 /* 0xec5c */;
                15128: data_o = 32'h00000000 /* 0xec60 */;
                15129: data_o = 32'h00000000 /* 0xec64 */;
                15130: data_o = 32'h00000000 /* 0xec68 */;
                15131: data_o = 32'h00000000 /* 0xec6c */;
                15132: data_o = 32'h00000000 /* 0xec70 */;
                15133: data_o = 32'h00000000 /* 0xec74 */;
                15134: data_o = 32'h00000000 /* 0xec78 */;
                15135: data_o = 32'h00000000 /* 0xec7c */;
                15136: data_o = 32'h00000000 /* 0xec80 */;
                15137: data_o = 32'h00000000 /* 0xec84 */;
                15138: data_o = 32'h00000000 /* 0xec88 */;
                15139: data_o = 32'h00000000 /* 0xec8c */;
                15140: data_o = 32'h00000000 /* 0xec90 */;
                15141: data_o = 32'h00000000 /* 0xec94 */;
                15142: data_o = 32'h00000000 /* 0xec98 */;
                15143: data_o = 32'h00000000 /* 0xec9c */;
                15144: data_o = 32'h00000000 /* 0xeca0 */;
                15145: data_o = 32'h00000000 /* 0xeca4 */;
                15146: data_o = 32'h00000000 /* 0xeca8 */;
                15147: data_o = 32'h00000000 /* 0xecac */;
                15148: data_o = 32'h00000000 /* 0xecb0 */;
                15149: data_o = 32'h00000000 /* 0xecb4 */;
                15150: data_o = 32'h00000000 /* 0xecb8 */;
                15151: data_o = 32'h00000000 /* 0xecbc */;
                15152: data_o = 32'h00000000 /* 0xecc0 */;
                15153: data_o = 32'h00000000 /* 0xecc4 */;
                15154: data_o = 32'h00000000 /* 0xecc8 */;
                15155: data_o = 32'h00000000 /* 0xeccc */;
                15156: data_o = 32'h00000000 /* 0xecd0 */;
                15157: data_o = 32'h00000000 /* 0xecd4 */;
                15158: data_o = 32'h00000000 /* 0xecd8 */;
                15159: data_o = 32'h00000000 /* 0xecdc */;
                15160: data_o = 32'h00000000 /* 0xece0 */;
                15161: data_o = 32'h00000000 /* 0xece4 */;
                15162: data_o = 32'h00000000 /* 0xece8 */;
                15163: data_o = 32'h00000000 /* 0xecec */;
                15164: data_o = 32'h00000000 /* 0xecf0 */;
                15165: data_o = 32'h00000000 /* 0xecf4 */;
                15166: data_o = 32'h00000000 /* 0xecf8 */;
                15167: data_o = 32'h00000000 /* 0xecfc */;
                15168: data_o = 32'h00000000 /* 0xed00 */;
                15169: data_o = 32'h00000000 /* 0xed04 */;
                15170: data_o = 32'h00000000 /* 0xed08 */;
                15171: data_o = 32'h00000000 /* 0xed0c */;
                15172: data_o = 32'h00000000 /* 0xed10 */;
                15173: data_o = 32'h00000000 /* 0xed14 */;
                15174: data_o = 32'h00000000 /* 0xed18 */;
                15175: data_o = 32'h00000000 /* 0xed1c */;
                15176: data_o = 32'h00000000 /* 0xed20 */;
                15177: data_o = 32'h00000000 /* 0xed24 */;
                15178: data_o = 32'h00000000 /* 0xed28 */;
                15179: data_o = 32'h00000000 /* 0xed2c */;
                15180: data_o = 32'h00000000 /* 0xed30 */;
                15181: data_o = 32'h00000000 /* 0xed34 */;
                15182: data_o = 32'h00000000 /* 0xed38 */;
                15183: data_o = 32'h00000000 /* 0xed3c */;
                15184: data_o = 32'h00000000 /* 0xed40 */;
                15185: data_o = 32'h00000000 /* 0xed44 */;
                15186: data_o = 32'h00000000 /* 0xed48 */;
                15187: data_o = 32'h00000000 /* 0xed4c */;
                15188: data_o = 32'h00000000 /* 0xed50 */;
                15189: data_o = 32'h00000000 /* 0xed54 */;
                15190: data_o = 32'h00000000 /* 0xed58 */;
                15191: data_o = 32'h00000000 /* 0xed5c */;
                15192: data_o = 32'h00000000 /* 0xed60 */;
                15193: data_o = 32'h00000000 /* 0xed64 */;
                15194: data_o = 32'h00000000 /* 0xed68 */;
                15195: data_o = 32'h00000000 /* 0xed6c */;
                15196: data_o = 32'h00000000 /* 0xed70 */;
                15197: data_o = 32'h00000000 /* 0xed74 */;
                15198: data_o = 32'h00000000 /* 0xed78 */;
                15199: data_o = 32'h00000000 /* 0xed7c */;
                15200: data_o = 32'h00000000 /* 0xed80 */;
                15201: data_o = 32'h00000000 /* 0xed84 */;
                15202: data_o = 32'h00000000 /* 0xed88 */;
                15203: data_o = 32'h00000000 /* 0xed8c */;
                15204: data_o = 32'h00000000 /* 0xed90 */;
                15205: data_o = 32'h00000000 /* 0xed94 */;
                15206: data_o = 32'h00000000 /* 0xed98 */;
                15207: data_o = 32'h00000000 /* 0xed9c */;
                15208: data_o = 32'h00000000 /* 0xeda0 */;
                15209: data_o = 32'h00000000 /* 0xeda4 */;
                15210: data_o = 32'h00000000 /* 0xeda8 */;
                15211: data_o = 32'h00000000 /* 0xedac */;
                15212: data_o = 32'h00000000 /* 0xedb0 */;
                15213: data_o = 32'h00000000 /* 0xedb4 */;
                15214: data_o = 32'h00000000 /* 0xedb8 */;
                15215: data_o = 32'h00000000 /* 0xedbc */;
                15216: data_o = 32'h00000000 /* 0xedc0 */;
                15217: data_o = 32'h00000000 /* 0xedc4 */;
                15218: data_o = 32'h00000000 /* 0xedc8 */;
                15219: data_o = 32'h00000000 /* 0xedcc */;
                15220: data_o = 32'h00000000 /* 0xedd0 */;
                15221: data_o = 32'h00000000 /* 0xedd4 */;
                15222: data_o = 32'h00000000 /* 0xedd8 */;
                15223: data_o = 32'h00000000 /* 0xeddc */;
                15224: data_o = 32'h00000000 /* 0xede0 */;
                15225: data_o = 32'h00000000 /* 0xede4 */;
                15226: data_o = 32'h00000000 /* 0xede8 */;
                15227: data_o = 32'h00000000 /* 0xedec */;
                15228: data_o = 32'h00000000 /* 0xedf0 */;
                15229: data_o = 32'h00000000 /* 0xedf4 */;
                15230: data_o = 32'h00000000 /* 0xedf8 */;
                15231: data_o = 32'h00000000 /* 0xedfc */;
                15232: data_o = 32'h00000000 /* 0xee00 */;
                15233: data_o = 32'h00000000 /* 0xee04 */;
                15234: data_o = 32'h00000000 /* 0xee08 */;
                15235: data_o = 32'h00000000 /* 0xee0c */;
                15236: data_o = 32'h00000000 /* 0xee10 */;
                15237: data_o = 32'h00000000 /* 0xee14 */;
                15238: data_o = 32'h00000000 /* 0xee18 */;
                15239: data_o = 32'h00000000 /* 0xee1c */;
                15240: data_o = 32'h00000000 /* 0xee20 */;
                15241: data_o = 32'h00000000 /* 0xee24 */;
                15242: data_o = 32'h00000000 /* 0xee28 */;
                15243: data_o = 32'h00000000 /* 0xee2c */;
                15244: data_o = 32'h00000000 /* 0xee30 */;
                15245: data_o = 32'h00000000 /* 0xee34 */;
                15246: data_o = 32'h00000000 /* 0xee38 */;
                15247: data_o = 32'h00000000 /* 0xee3c */;
                15248: data_o = 32'h00000000 /* 0xee40 */;
                15249: data_o = 32'h00000000 /* 0xee44 */;
                15250: data_o = 32'h00000000 /* 0xee48 */;
                15251: data_o = 32'h00000000 /* 0xee4c */;
                15252: data_o = 32'h00000000 /* 0xee50 */;
                15253: data_o = 32'h00000000 /* 0xee54 */;
                15254: data_o = 32'h00000000 /* 0xee58 */;
                15255: data_o = 32'h00000000 /* 0xee5c */;
                15256: data_o = 32'h00000000 /* 0xee60 */;
                15257: data_o = 32'h00000000 /* 0xee64 */;
                15258: data_o = 32'h00000000 /* 0xee68 */;
                15259: data_o = 32'h00000000 /* 0xee6c */;
                15260: data_o = 32'h00000000 /* 0xee70 */;
                15261: data_o = 32'h00000000 /* 0xee74 */;
                15262: data_o = 32'h00000000 /* 0xee78 */;
                15263: data_o = 32'h00000000 /* 0xee7c */;
                15264: data_o = 32'h00000000 /* 0xee80 */;
                15265: data_o = 32'h00000000 /* 0xee84 */;
                15266: data_o = 32'h00000000 /* 0xee88 */;
                15267: data_o = 32'h00000000 /* 0xee8c */;
                15268: data_o = 32'h00000000 /* 0xee90 */;
                15269: data_o = 32'h00000000 /* 0xee94 */;
                15270: data_o = 32'h00000000 /* 0xee98 */;
                15271: data_o = 32'h00000000 /* 0xee9c */;
                15272: data_o = 32'h00000000 /* 0xeea0 */;
                15273: data_o = 32'h00000000 /* 0xeea4 */;
                15274: data_o = 32'h00000000 /* 0xeea8 */;
                15275: data_o = 32'h00000000 /* 0xeeac */;
                15276: data_o = 32'h00000000 /* 0xeeb0 */;
                15277: data_o = 32'h00000000 /* 0xeeb4 */;
                15278: data_o = 32'h00000000 /* 0xeeb8 */;
                15279: data_o = 32'h00000000 /* 0xeebc */;
                15280: data_o = 32'h00000000 /* 0xeec0 */;
                15281: data_o = 32'h00000000 /* 0xeec4 */;
                15282: data_o = 32'h00000000 /* 0xeec8 */;
                15283: data_o = 32'h00000000 /* 0xeecc */;
                15284: data_o = 32'h00000000 /* 0xeed0 */;
                15285: data_o = 32'h00000000 /* 0xeed4 */;
                15286: data_o = 32'h00000000 /* 0xeed8 */;
                15287: data_o = 32'h00000000 /* 0xeedc */;
                15288: data_o = 32'h00000000 /* 0xeee0 */;
                15289: data_o = 32'h00000000 /* 0xeee4 */;
                15290: data_o = 32'h00000000 /* 0xeee8 */;
                15291: data_o = 32'h00000000 /* 0xeeec */;
                15292: data_o = 32'h00000000 /* 0xeef0 */;
                15293: data_o = 32'h00000000 /* 0xeef4 */;
                15294: data_o = 32'h00000000 /* 0xeef8 */;
                15295: data_o = 32'h00000000 /* 0xeefc */;
                15296: data_o = 32'h00000000 /* 0xef00 */;
                15297: data_o = 32'h00000000 /* 0xef04 */;
                15298: data_o = 32'h00000000 /* 0xef08 */;
                15299: data_o = 32'h00000000 /* 0xef0c */;
                15300: data_o = 32'h00000000 /* 0xef10 */;
                15301: data_o = 32'h00000000 /* 0xef14 */;
                15302: data_o = 32'h00000000 /* 0xef18 */;
                15303: data_o = 32'h00000000 /* 0xef1c */;
                15304: data_o = 32'h00000000 /* 0xef20 */;
                15305: data_o = 32'h00000000 /* 0xef24 */;
                15306: data_o = 32'h00000000 /* 0xef28 */;
                15307: data_o = 32'h00000000 /* 0xef2c */;
                15308: data_o = 32'h00000000 /* 0xef30 */;
                15309: data_o = 32'h00000000 /* 0xef34 */;
                15310: data_o = 32'h00000000 /* 0xef38 */;
                15311: data_o = 32'h00000000 /* 0xef3c */;
                15312: data_o = 32'h00000000 /* 0xef40 */;
                15313: data_o = 32'h00000000 /* 0xef44 */;
                15314: data_o = 32'h00000000 /* 0xef48 */;
                15315: data_o = 32'h00000000 /* 0xef4c */;
                15316: data_o = 32'h00000000 /* 0xef50 */;
                15317: data_o = 32'h00000000 /* 0xef54 */;
                15318: data_o = 32'h00000000 /* 0xef58 */;
                15319: data_o = 32'h00000000 /* 0xef5c */;
                15320: data_o = 32'h00000000 /* 0xef60 */;
                15321: data_o = 32'h00000000 /* 0xef64 */;
                15322: data_o = 32'h00000000 /* 0xef68 */;
                15323: data_o = 32'h00000000 /* 0xef6c */;
                15324: data_o = 32'h00000000 /* 0xef70 */;
                15325: data_o = 32'h00000000 /* 0xef74 */;
                15326: data_o = 32'h00000000 /* 0xef78 */;
                15327: data_o = 32'h00000000 /* 0xef7c */;
                15328: data_o = 32'h00000000 /* 0xef80 */;
                15329: data_o = 32'h00000000 /* 0xef84 */;
                15330: data_o = 32'h00000000 /* 0xef88 */;
                15331: data_o = 32'h00000000 /* 0xef8c */;
                15332: data_o = 32'h00000000 /* 0xef90 */;
                15333: data_o = 32'h00000000 /* 0xef94 */;
                15334: data_o = 32'h00000000 /* 0xef98 */;
                15335: data_o = 32'h00000000 /* 0xef9c */;
                15336: data_o = 32'h00000000 /* 0xefa0 */;
                15337: data_o = 32'h00000000 /* 0xefa4 */;
                15338: data_o = 32'h00000000 /* 0xefa8 */;
                15339: data_o = 32'h00000000 /* 0xefac */;
                15340: data_o = 32'h00000000 /* 0xefb0 */;
                15341: data_o = 32'h00000000 /* 0xefb4 */;
                15342: data_o = 32'h00000000 /* 0xefb8 */;
                15343: data_o = 32'h00000000 /* 0xefbc */;
                15344: data_o = 32'h00000000 /* 0xefc0 */;
                15345: data_o = 32'h00000000 /* 0xefc4 */;
                15346: data_o = 32'h00000000 /* 0xefc8 */;
                15347: data_o = 32'h00000000 /* 0xefcc */;
                15348: data_o = 32'h00000000 /* 0xefd0 */;
                15349: data_o = 32'h00000000 /* 0xefd4 */;
                15350: data_o = 32'h00000000 /* 0xefd8 */;
                15351: data_o = 32'h00000000 /* 0xefdc */;
                15352: data_o = 32'h00000000 /* 0xefe0 */;
                15353: data_o = 32'h00000000 /* 0xefe4 */;
                15354: data_o = 32'h00000000 /* 0xefe8 */;
                15355: data_o = 32'h00000000 /* 0xefec */;
                15356: data_o = 32'h00000000 /* 0xeff0 */;
                15357: data_o = 32'h00000000 /* 0xeff4 */;
                15358: data_o = 32'h00000000 /* 0xeff8 */;
                15359: data_o = 32'h00000000 /* 0xeffc */;
                15360: data_o = 32'h00000000 /* 0xf000 */;
                15361: data_o = 32'h00000000 /* 0xf004 */;
                15362: data_o = 32'h00000000 /* 0xf008 */;
                15363: data_o = 32'h00000000 /* 0xf00c */;
                15364: data_o = 32'h00000000 /* 0xf010 */;
                15365: data_o = 32'h00000000 /* 0xf014 */;
                15366: data_o = 32'h00000000 /* 0xf018 */;
                15367: data_o = 32'h00000000 /* 0xf01c */;
                15368: data_o = 32'h00000000 /* 0xf020 */;
                15369: data_o = 32'h00000000 /* 0xf024 */;
                15370: data_o = 32'h00000000 /* 0xf028 */;
                15371: data_o = 32'h00000000 /* 0xf02c */;
                15372: data_o = 32'h00000000 /* 0xf030 */;
                15373: data_o = 32'h00000000 /* 0xf034 */;
                15374: data_o = 32'h00000000 /* 0xf038 */;
                15375: data_o = 32'h00000000 /* 0xf03c */;
                15376: data_o = 32'h00000000 /* 0xf040 */;
                15377: data_o = 32'h00000000 /* 0xf044 */;
                15378: data_o = 32'h00000000 /* 0xf048 */;
                15379: data_o = 32'h00000000 /* 0xf04c */;
                15380: data_o = 32'h00000000 /* 0xf050 */;
                15381: data_o = 32'h00000000 /* 0xf054 */;
                15382: data_o = 32'h00000000 /* 0xf058 */;
                15383: data_o = 32'h00000000 /* 0xf05c */;
                15384: data_o = 32'h00000000 /* 0xf060 */;
                15385: data_o = 32'h00000000 /* 0xf064 */;
                15386: data_o = 32'h00000000 /* 0xf068 */;
                15387: data_o = 32'h00000000 /* 0xf06c */;
                15388: data_o = 32'h00000000 /* 0xf070 */;
                15389: data_o = 32'h00000000 /* 0xf074 */;
                15390: data_o = 32'h00000000 /* 0xf078 */;
                15391: data_o = 32'h00000000 /* 0xf07c */;
                15392: data_o = 32'h00000000 /* 0xf080 */;
                15393: data_o = 32'h00000000 /* 0xf084 */;
                15394: data_o = 32'h00000000 /* 0xf088 */;
                15395: data_o = 32'h00000000 /* 0xf08c */;
                15396: data_o = 32'h00000000 /* 0xf090 */;
                15397: data_o = 32'h00000000 /* 0xf094 */;
                15398: data_o = 32'h00000000 /* 0xf098 */;
                15399: data_o = 32'h00000000 /* 0xf09c */;
                15400: data_o = 32'h00000000 /* 0xf0a0 */;
                15401: data_o = 32'h00000000 /* 0xf0a4 */;
                15402: data_o = 32'h00000000 /* 0xf0a8 */;
                15403: data_o = 32'h00000000 /* 0xf0ac */;
                15404: data_o = 32'h00000000 /* 0xf0b0 */;
                15405: data_o = 32'h00000000 /* 0xf0b4 */;
                15406: data_o = 32'h00000000 /* 0xf0b8 */;
                15407: data_o = 32'h00000000 /* 0xf0bc */;
                15408: data_o = 32'h00000000 /* 0xf0c0 */;
                15409: data_o = 32'h00000000 /* 0xf0c4 */;
                15410: data_o = 32'h00000000 /* 0xf0c8 */;
                15411: data_o = 32'h00000000 /* 0xf0cc */;
                15412: data_o = 32'h00000000 /* 0xf0d0 */;
                15413: data_o = 32'h00000000 /* 0xf0d4 */;
                15414: data_o = 32'h00000000 /* 0xf0d8 */;
                15415: data_o = 32'h00000000 /* 0xf0dc */;
                15416: data_o = 32'h00000000 /* 0xf0e0 */;
                15417: data_o = 32'h00000000 /* 0xf0e4 */;
                15418: data_o = 32'h00000000 /* 0xf0e8 */;
                15419: data_o = 32'h00000000 /* 0xf0ec */;
                15420: data_o = 32'h00000000 /* 0xf0f0 */;
                15421: data_o = 32'h00000000 /* 0xf0f4 */;
                15422: data_o = 32'h00000000 /* 0xf0f8 */;
                15423: data_o = 32'h00000000 /* 0xf0fc */;
                15424: data_o = 32'h00000000 /* 0xf100 */;
                15425: data_o = 32'h00000000 /* 0xf104 */;
                15426: data_o = 32'h00000000 /* 0xf108 */;
                15427: data_o = 32'h00000000 /* 0xf10c */;
                15428: data_o = 32'h00000000 /* 0xf110 */;
                15429: data_o = 32'h00000000 /* 0xf114 */;
                15430: data_o = 32'h00000000 /* 0xf118 */;
                15431: data_o = 32'h00000000 /* 0xf11c */;
                15432: data_o = 32'h00000000 /* 0xf120 */;
                15433: data_o = 32'h00000000 /* 0xf124 */;
                15434: data_o = 32'h00000000 /* 0xf128 */;
                15435: data_o = 32'h00000000 /* 0xf12c */;
                15436: data_o = 32'h00000000 /* 0xf130 */;
                15437: data_o = 32'h00000000 /* 0xf134 */;
                15438: data_o = 32'h00000000 /* 0xf138 */;
                15439: data_o = 32'h00000000 /* 0xf13c */;
                15440: data_o = 32'h00000000 /* 0xf140 */;
                15441: data_o = 32'h00000000 /* 0xf144 */;
                15442: data_o = 32'h00000000 /* 0xf148 */;
                15443: data_o = 32'h00000000 /* 0xf14c */;
                15444: data_o = 32'h00000000 /* 0xf150 */;
                15445: data_o = 32'h00000000 /* 0xf154 */;
                15446: data_o = 32'h00000000 /* 0xf158 */;
                15447: data_o = 32'h00000000 /* 0xf15c */;
                15448: data_o = 32'h00000000 /* 0xf160 */;
                15449: data_o = 32'h00000000 /* 0xf164 */;
                15450: data_o = 32'h00000000 /* 0xf168 */;
                15451: data_o = 32'h00000000 /* 0xf16c */;
                15452: data_o = 32'h00000000 /* 0xf170 */;
                15453: data_o = 32'h00000000 /* 0xf174 */;
                15454: data_o = 32'h00000000 /* 0xf178 */;
                15455: data_o = 32'h00000000 /* 0xf17c */;
                15456: data_o = 32'h00000000 /* 0xf180 */;
                15457: data_o = 32'h00000000 /* 0xf184 */;
                15458: data_o = 32'h00000000 /* 0xf188 */;
                15459: data_o = 32'h00000000 /* 0xf18c */;
                15460: data_o = 32'h00000000 /* 0xf190 */;
                15461: data_o = 32'h00000000 /* 0xf194 */;
                15462: data_o = 32'h00000000 /* 0xf198 */;
                15463: data_o = 32'h00000000 /* 0xf19c */;
                15464: data_o = 32'h00000000 /* 0xf1a0 */;
                15465: data_o = 32'h00000000 /* 0xf1a4 */;
                15466: data_o = 32'h00000000 /* 0xf1a8 */;
                15467: data_o = 32'h00000000 /* 0xf1ac */;
                15468: data_o = 32'h00000000 /* 0xf1b0 */;
                15469: data_o = 32'h00000000 /* 0xf1b4 */;
                15470: data_o = 32'h00000000 /* 0xf1b8 */;
                15471: data_o = 32'h00000000 /* 0xf1bc */;
                15472: data_o = 32'h00000000 /* 0xf1c0 */;
                15473: data_o = 32'h00000000 /* 0xf1c4 */;
                15474: data_o = 32'h00000000 /* 0xf1c8 */;
                15475: data_o = 32'h00000000 /* 0xf1cc */;
                15476: data_o = 32'h00000000 /* 0xf1d0 */;
                15477: data_o = 32'h00000000 /* 0xf1d4 */;
                15478: data_o = 32'h00000000 /* 0xf1d8 */;
                15479: data_o = 32'h00000000 /* 0xf1dc */;
                15480: data_o = 32'h00000000 /* 0xf1e0 */;
                15481: data_o = 32'h00000000 /* 0xf1e4 */;
                15482: data_o = 32'h00000000 /* 0xf1e8 */;
                15483: data_o = 32'h00000000 /* 0xf1ec */;
                15484: data_o = 32'h00000000 /* 0xf1f0 */;
                15485: data_o = 32'h00000000 /* 0xf1f4 */;
                15486: data_o = 32'h00000000 /* 0xf1f8 */;
                15487: data_o = 32'h00000000 /* 0xf1fc */;
                15488: data_o = 32'h00000000 /* 0xf200 */;
                15489: data_o = 32'h00000000 /* 0xf204 */;
                15490: data_o = 32'h00000000 /* 0xf208 */;
                15491: data_o = 32'h00000000 /* 0xf20c */;
                15492: data_o = 32'h00000000 /* 0xf210 */;
                15493: data_o = 32'h00000000 /* 0xf214 */;
                15494: data_o = 32'h00000000 /* 0xf218 */;
                15495: data_o = 32'h00000000 /* 0xf21c */;
                15496: data_o = 32'h00000000 /* 0xf220 */;
                15497: data_o = 32'h00000000 /* 0xf224 */;
                15498: data_o = 32'h00000000 /* 0xf228 */;
                15499: data_o = 32'h00000000 /* 0xf22c */;
                15500: data_o = 32'h00000000 /* 0xf230 */;
                15501: data_o = 32'h00000000 /* 0xf234 */;
                15502: data_o = 32'h00000000 /* 0xf238 */;
                15503: data_o = 32'h00000000 /* 0xf23c */;
                15504: data_o = 32'h00000000 /* 0xf240 */;
                15505: data_o = 32'h00000000 /* 0xf244 */;
                15506: data_o = 32'h00000000 /* 0xf248 */;
                15507: data_o = 32'h00000000 /* 0xf24c */;
                15508: data_o = 32'h00000000 /* 0xf250 */;
                15509: data_o = 32'h00000000 /* 0xf254 */;
                15510: data_o = 32'h00000000 /* 0xf258 */;
                15511: data_o = 32'h00000000 /* 0xf25c */;
                15512: data_o = 32'h00000000 /* 0xf260 */;
                15513: data_o = 32'h00000000 /* 0xf264 */;
                15514: data_o = 32'h00000000 /* 0xf268 */;
                15515: data_o = 32'h00000000 /* 0xf26c */;
                15516: data_o = 32'h00000000 /* 0xf270 */;
                15517: data_o = 32'h00000000 /* 0xf274 */;
                15518: data_o = 32'h00000000 /* 0xf278 */;
                15519: data_o = 32'h00000000 /* 0xf27c */;
                15520: data_o = 32'h00000000 /* 0xf280 */;
                15521: data_o = 32'h00000000 /* 0xf284 */;
                15522: data_o = 32'h00000000 /* 0xf288 */;
                15523: data_o = 32'h00000000 /* 0xf28c */;
                15524: data_o = 32'h00000000 /* 0xf290 */;
                15525: data_o = 32'h00000000 /* 0xf294 */;
                15526: data_o = 32'h00000000 /* 0xf298 */;
                15527: data_o = 32'h00000000 /* 0xf29c */;
                15528: data_o = 32'h00000000 /* 0xf2a0 */;
                15529: data_o = 32'h00000000 /* 0xf2a4 */;
                15530: data_o = 32'h00000000 /* 0xf2a8 */;
                15531: data_o = 32'h00000000 /* 0xf2ac */;
                15532: data_o = 32'h00000000 /* 0xf2b0 */;
                15533: data_o = 32'h00000000 /* 0xf2b4 */;
                15534: data_o = 32'h00000000 /* 0xf2b8 */;
                15535: data_o = 32'h00000000 /* 0xf2bc */;
                15536: data_o = 32'h00000000 /* 0xf2c0 */;
                15537: data_o = 32'h00000000 /* 0xf2c4 */;
                15538: data_o = 32'h00000000 /* 0xf2c8 */;
                15539: data_o = 32'h00000000 /* 0xf2cc */;
                15540: data_o = 32'h00000000 /* 0xf2d0 */;
                15541: data_o = 32'h00000000 /* 0xf2d4 */;
                15542: data_o = 32'h00000000 /* 0xf2d8 */;
                15543: data_o = 32'h00000000 /* 0xf2dc */;
                15544: data_o = 32'h00000000 /* 0xf2e0 */;
                15545: data_o = 32'h00000000 /* 0xf2e4 */;
                15546: data_o = 32'h00000000 /* 0xf2e8 */;
                15547: data_o = 32'h00000000 /* 0xf2ec */;
                15548: data_o = 32'h00000000 /* 0xf2f0 */;
                15549: data_o = 32'h00000000 /* 0xf2f4 */;
                15550: data_o = 32'h00000000 /* 0xf2f8 */;
                15551: data_o = 32'h00000000 /* 0xf2fc */;
                15552: data_o = 32'h00000000 /* 0xf300 */;
                15553: data_o = 32'h00000000 /* 0xf304 */;
                15554: data_o = 32'h00000000 /* 0xf308 */;
                15555: data_o = 32'h00000000 /* 0xf30c */;
                15556: data_o = 32'h00000000 /* 0xf310 */;
                15557: data_o = 32'h00000000 /* 0xf314 */;
                15558: data_o = 32'h00000000 /* 0xf318 */;
                15559: data_o = 32'h00000000 /* 0xf31c */;
                15560: data_o = 32'h00000000 /* 0xf320 */;
                15561: data_o = 32'h00000000 /* 0xf324 */;
                15562: data_o = 32'h00000000 /* 0xf328 */;
                15563: data_o = 32'h00000000 /* 0xf32c */;
                15564: data_o = 32'h00000000 /* 0xf330 */;
                15565: data_o = 32'h00000000 /* 0xf334 */;
                15566: data_o = 32'h00000000 /* 0xf338 */;
                15567: data_o = 32'h00000000 /* 0xf33c */;
                15568: data_o = 32'h00000000 /* 0xf340 */;
                15569: data_o = 32'h00000000 /* 0xf344 */;
                15570: data_o = 32'h00000000 /* 0xf348 */;
                15571: data_o = 32'h00000000 /* 0xf34c */;
                15572: data_o = 32'h00000000 /* 0xf350 */;
                15573: data_o = 32'h00000000 /* 0xf354 */;
                15574: data_o = 32'h00000000 /* 0xf358 */;
                15575: data_o = 32'h00000000 /* 0xf35c */;
                15576: data_o = 32'h00000000 /* 0xf360 */;
                15577: data_o = 32'h00000000 /* 0xf364 */;
                15578: data_o = 32'h00000000 /* 0xf368 */;
                15579: data_o = 32'h00000000 /* 0xf36c */;
                15580: data_o = 32'h00000000 /* 0xf370 */;
                15581: data_o = 32'h00000000 /* 0xf374 */;
                15582: data_o = 32'h00000000 /* 0xf378 */;
                15583: data_o = 32'h00000000 /* 0xf37c */;
                15584: data_o = 32'h00000000 /* 0xf380 */;
                15585: data_o = 32'h00000000 /* 0xf384 */;
                15586: data_o = 32'h00000000 /* 0xf388 */;
                15587: data_o = 32'h00000000 /* 0xf38c */;
                15588: data_o = 32'h00000000 /* 0xf390 */;
                15589: data_o = 32'h00000000 /* 0xf394 */;
                15590: data_o = 32'h00000000 /* 0xf398 */;
                15591: data_o = 32'h00000000 /* 0xf39c */;
                15592: data_o = 32'h00000000 /* 0xf3a0 */;
                15593: data_o = 32'h00000000 /* 0xf3a4 */;
                15594: data_o = 32'h00000000 /* 0xf3a8 */;
                15595: data_o = 32'h00000000 /* 0xf3ac */;
                15596: data_o = 32'h00000000 /* 0xf3b0 */;
                15597: data_o = 32'h00000000 /* 0xf3b4 */;
                15598: data_o = 32'h00000000 /* 0xf3b8 */;
                15599: data_o = 32'h00000000 /* 0xf3bc */;
                15600: data_o = 32'h00000000 /* 0xf3c0 */;
                15601: data_o = 32'h00000000 /* 0xf3c4 */;
                15602: data_o = 32'h00000000 /* 0xf3c8 */;
                15603: data_o = 32'h00000000 /* 0xf3cc */;
                15604: data_o = 32'h00000000 /* 0xf3d0 */;
                15605: data_o = 32'h00000000 /* 0xf3d4 */;
                15606: data_o = 32'h00000000 /* 0xf3d8 */;
                15607: data_o = 32'h00000000 /* 0xf3dc */;
                15608: data_o = 32'h00000000 /* 0xf3e0 */;
                15609: data_o = 32'h00000000 /* 0xf3e4 */;
                15610: data_o = 32'h00000000 /* 0xf3e8 */;
                15611: data_o = 32'h00000000 /* 0xf3ec */;
                15612: data_o = 32'h00000000 /* 0xf3f0 */;
                15613: data_o = 32'h00000000 /* 0xf3f4 */;
                15614: data_o = 32'h00000000 /* 0xf3f8 */;
                15615: data_o = 32'h00000000 /* 0xf3fc */;
                15616: data_o = 32'h00000000 /* 0xf400 */;
                15617: data_o = 32'h00000000 /* 0xf404 */;
                15618: data_o = 32'h00000000 /* 0xf408 */;
                15619: data_o = 32'h00000000 /* 0xf40c */;
                15620: data_o = 32'h00000000 /* 0xf410 */;
                15621: data_o = 32'h00000000 /* 0xf414 */;
                15622: data_o = 32'h00000000 /* 0xf418 */;
                15623: data_o = 32'h00000000 /* 0xf41c */;
                15624: data_o = 32'h00000000 /* 0xf420 */;
                15625: data_o = 32'h00000000 /* 0xf424 */;
                15626: data_o = 32'h00000000 /* 0xf428 */;
                15627: data_o = 32'h00000000 /* 0xf42c */;
                15628: data_o = 32'h00000000 /* 0xf430 */;
                15629: data_o = 32'h00000000 /* 0xf434 */;
                15630: data_o = 32'h00000000 /* 0xf438 */;
                15631: data_o = 32'h00000000 /* 0xf43c */;
                15632: data_o = 32'h00000000 /* 0xf440 */;
                15633: data_o = 32'h00000000 /* 0xf444 */;
                15634: data_o = 32'h00000000 /* 0xf448 */;
                15635: data_o = 32'h00000000 /* 0xf44c */;
                15636: data_o = 32'h00000000 /* 0xf450 */;
                15637: data_o = 32'h00000000 /* 0xf454 */;
                15638: data_o = 32'h00000000 /* 0xf458 */;
                15639: data_o = 32'h00000000 /* 0xf45c */;
                15640: data_o = 32'h00000000 /* 0xf460 */;
                15641: data_o = 32'h00000000 /* 0xf464 */;
                15642: data_o = 32'h00000000 /* 0xf468 */;
                15643: data_o = 32'h00000000 /* 0xf46c */;
                15644: data_o = 32'h00000000 /* 0xf470 */;
                15645: data_o = 32'h00000000 /* 0xf474 */;
                15646: data_o = 32'h00000000 /* 0xf478 */;
                15647: data_o = 32'h00000000 /* 0xf47c */;
                15648: data_o = 32'h00000000 /* 0xf480 */;
                15649: data_o = 32'h00000000 /* 0xf484 */;
                15650: data_o = 32'h00000000 /* 0xf488 */;
                15651: data_o = 32'h00000000 /* 0xf48c */;
                15652: data_o = 32'h00000000 /* 0xf490 */;
                15653: data_o = 32'h00000000 /* 0xf494 */;
                15654: data_o = 32'h00000000 /* 0xf498 */;
                15655: data_o = 32'h00000000 /* 0xf49c */;
                15656: data_o = 32'h00000000 /* 0xf4a0 */;
                15657: data_o = 32'h00000000 /* 0xf4a4 */;
                15658: data_o = 32'h00000000 /* 0xf4a8 */;
                15659: data_o = 32'h00000000 /* 0xf4ac */;
                15660: data_o = 32'h00000000 /* 0xf4b0 */;
                15661: data_o = 32'h00000000 /* 0xf4b4 */;
                15662: data_o = 32'h00000000 /* 0xf4b8 */;
                15663: data_o = 32'h00000000 /* 0xf4bc */;
                15664: data_o = 32'h00000000 /* 0xf4c0 */;
                15665: data_o = 32'h00000000 /* 0xf4c4 */;
                15666: data_o = 32'h00000000 /* 0xf4c8 */;
                15667: data_o = 32'h00000000 /* 0xf4cc */;
                15668: data_o = 32'h00000000 /* 0xf4d0 */;
                15669: data_o = 32'h00000000 /* 0xf4d4 */;
                15670: data_o = 32'h00000000 /* 0xf4d8 */;
                15671: data_o = 32'h00000000 /* 0xf4dc */;
                15672: data_o = 32'h00000000 /* 0xf4e0 */;
                15673: data_o = 32'h00000000 /* 0xf4e4 */;
                15674: data_o = 32'h00000000 /* 0xf4e8 */;
                15675: data_o = 32'h00000000 /* 0xf4ec */;
                15676: data_o = 32'h00000000 /* 0xf4f0 */;
                15677: data_o = 32'h00000000 /* 0xf4f4 */;
                15678: data_o = 32'h00000000 /* 0xf4f8 */;
                15679: data_o = 32'h00000000 /* 0xf4fc */;
                15680: data_o = 32'h00000000 /* 0xf500 */;
                15681: data_o = 32'h00000000 /* 0xf504 */;
                15682: data_o = 32'h00000000 /* 0xf508 */;
                15683: data_o = 32'h00000000 /* 0xf50c */;
                15684: data_o = 32'h00000000 /* 0xf510 */;
                15685: data_o = 32'h00000000 /* 0xf514 */;
                15686: data_o = 32'h00000000 /* 0xf518 */;
                15687: data_o = 32'h00000000 /* 0xf51c */;
                15688: data_o = 32'h00000000 /* 0xf520 */;
                15689: data_o = 32'h00000000 /* 0xf524 */;
                15690: data_o = 32'h00000000 /* 0xf528 */;
                15691: data_o = 32'h00000000 /* 0xf52c */;
                15692: data_o = 32'h00000000 /* 0xf530 */;
                15693: data_o = 32'h00000000 /* 0xf534 */;
                15694: data_o = 32'h00000000 /* 0xf538 */;
                15695: data_o = 32'h00000000 /* 0xf53c */;
                15696: data_o = 32'h00000000 /* 0xf540 */;
                15697: data_o = 32'h00000000 /* 0xf544 */;
                15698: data_o = 32'h00000000 /* 0xf548 */;
                15699: data_o = 32'h00000000 /* 0xf54c */;
                15700: data_o = 32'h00000000 /* 0xf550 */;
                15701: data_o = 32'h00000000 /* 0xf554 */;
                15702: data_o = 32'h00000000 /* 0xf558 */;
                15703: data_o = 32'h00000000 /* 0xf55c */;
                15704: data_o = 32'h00000000 /* 0xf560 */;
                15705: data_o = 32'h00000000 /* 0xf564 */;
                15706: data_o = 32'h00000000 /* 0xf568 */;
                15707: data_o = 32'h00000000 /* 0xf56c */;
                15708: data_o = 32'h00000000 /* 0xf570 */;
                15709: data_o = 32'h00000000 /* 0xf574 */;
                15710: data_o = 32'h00000000 /* 0xf578 */;
                15711: data_o = 32'h00000000 /* 0xf57c */;
                15712: data_o = 32'h00000000 /* 0xf580 */;
                15713: data_o = 32'h00000000 /* 0xf584 */;
                15714: data_o = 32'h00000000 /* 0xf588 */;
                15715: data_o = 32'h00000000 /* 0xf58c */;
                15716: data_o = 32'h00000000 /* 0xf590 */;
                15717: data_o = 32'h00000000 /* 0xf594 */;
                15718: data_o = 32'h00000000 /* 0xf598 */;
                15719: data_o = 32'h00000000 /* 0xf59c */;
                15720: data_o = 32'h00000000 /* 0xf5a0 */;
                15721: data_o = 32'h00000000 /* 0xf5a4 */;
                15722: data_o = 32'h00000000 /* 0xf5a8 */;
                15723: data_o = 32'h00000000 /* 0xf5ac */;
                15724: data_o = 32'h00000000 /* 0xf5b0 */;
                15725: data_o = 32'h00000000 /* 0xf5b4 */;
                15726: data_o = 32'h00000000 /* 0xf5b8 */;
                15727: data_o = 32'h00000000 /* 0xf5bc */;
                15728: data_o = 32'h00000000 /* 0xf5c0 */;
                15729: data_o = 32'h00000000 /* 0xf5c4 */;
                15730: data_o = 32'h00000000 /* 0xf5c8 */;
                15731: data_o = 32'h00000000 /* 0xf5cc */;
                15732: data_o = 32'h00000000 /* 0xf5d0 */;
                15733: data_o = 32'h00000000 /* 0xf5d4 */;
                15734: data_o = 32'h00000000 /* 0xf5d8 */;
                15735: data_o = 32'h00000000 /* 0xf5dc */;
                15736: data_o = 32'h00000000 /* 0xf5e0 */;
                15737: data_o = 32'h00000000 /* 0xf5e4 */;
                15738: data_o = 32'h00000000 /* 0xf5e8 */;
                15739: data_o = 32'h00000000 /* 0xf5ec */;
                15740: data_o = 32'h00000000 /* 0xf5f0 */;
                15741: data_o = 32'h00000000 /* 0xf5f4 */;
                15742: data_o = 32'h00000000 /* 0xf5f8 */;
                15743: data_o = 32'h00000000 /* 0xf5fc */;
                15744: data_o = 32'h00000000 /* 0xf600 */;
                15745: data_o = 32'h00000000 /* 0xf604 */;
                15746: data_o = 32'h00000000 /* 0xf608 */;
                15747: data_o = 32'h00000000 /* 0xf60c */;
                15748: data_o = 32'h00000000 /* 0xf610 */;
                15749: data_o = 32'h00000000 /* 0xf614 */;
                15750: data_o = 32'h00000000 /* 0xf618 */;
                15751: data_o = 32'h00000000 /* 0xf61c */;
                15752: data_o = 32'h00000000 /* 0xf620 */;
                15753: data_o = 32'h00000000 /* 0xf624 */;
                15754: data_o = 32'h00000000 /* 0xf628 */;
                15755: data_o = 32'h00000000 /* 0xf62c */;
                15756: data_o = 32'h00000000 /* 0xf630 */;
                15757: data_o = 32'h00000000 /* 0xf634 */;
                15758: data_o = 32'h00000000 /* 0xf638 */;
                15759: data_o = 32'h00000000 /* 0xf63c */;
                15760: data_o = 32'h00000000 /* 0xf640 */;
                15761: data_o = 32'h00000000 /* 0xf644 */;
                15762: data_o = 32'h00000000 /* 0xf648 */;
                15763: data_o = 32'h00000000 /* 0xf64c */;
                15764: data_o = 32'h00000000 /* 0xf650 */;
                15765: data_o = 32'h00000000 /* 0xf654 */;
                15766: data_o = 32'h00000000 /* 0xf658 */;
                15767: data_o = 32'h00000000 /* 0xf65c */;
                15768: data_o = 32'h00000000 /* 0xf660 */;
                15769: data_o = 32'h00000000 /* 0xf664 */;
                15770: data_o = 32'h00000000 /* 0xf668 */;
                15771: data_o = 32'h00000000 /* 0xf66c */;
                15772: data_o = 32'h00000000 /* 0xf670 */;
                15773: data_o = 32'h00000000 /* 0xf674 */;
                15774: data_o = 32'h00000000 /* 0xf678 */;
                15775: data_o = 32'h00000000 /* 0xf67c */;
                15776: data_o = 32'h00000000 /* 0xf680 */;
                15777: data_o = 32'h00000000 /* 0xf684 */;
                15778: data_o = 32'h00000000 /* 0xf688 */;
                15779: data_o = 32'h00000000 /* 0xf68c */;
                15780: data_o = 32'h00000000 /* 0xf690 */;
                15781: data_o = 32'h00000000 /* 0xf694 */;
                15782: data_o = 32'h00000000 /* 0xf698 */;
                15783: data_o = 32'h00000000 /* 0xf69c */;
                15784: data_o = 32'h00000000 /* 0xf6a0 */;
                15785: data_o = 32'h00000000 /* 0xf6a4 */;
                15786: data_o = 32'h00000000 /* 0xf6a8 */;
                15787: data_o = 32'h00000000 /* 0xf6ac */;
                15788: data_o = 32'h00000000 /* 0xf6b0 */;
                15789: data_o = 32'h00000000 /* 0xf6b4 */;
                15790: data_o = 32'h00000000 /* 0xf6b8 */;
                15791: data_o = 32'h00000000 /* 0xf6bc */;
                15792: data_o = 32'h00000000 /* 0xf6c0 */;
                15793: data_o = 32'h00000000 /* 0xf6c4 */;
                15794: data_o = 32'h00000000 /* 0xf6c8 */;
                15795: data_o = 32'h00000000 /* 0xf6cc */;
                15796: data_o = 32'h00000000 /* 0xf6d0 */;
                15797: data_o = 32'h00000000 /* 0xf6d4 */;
                15798: data_o = 32'h00000000 /* 0xf6d8 */;
                15799: data_o = 32'h00000000 /* 0xf6dc */;
                15800: data_o = 32'h00000000 /* 0xf6e0 */;
                15801: data_o = 32'h00000000 /* 0xf6e4 */;
                15802: data_o = 32'h00000000 /* 0xf6e8 */;
                15803: data_o = 32'h00000000 /* 0xf6ec */;
                15804: data_o = 32'h00000000 /* 0xf6f0 */;
                15805: data_o = 32'h00000000 /* 0xf6f4 */;
                15806: data_o = 32'h00000000 /* 0xf6f8 */;
                15807: data_o = 32'h00000000 /* 0xf6fc */;
                15808: data_o = 32'h00000000 /* 0xf700 */;
                15809: data_o = 32'h00000000 /* 0xf704 */;
                15810: data_o = 32'h00000000 /* 0xf708 */;
                15811: data_o = 32'h00000000 /* 0xf70c */;
                15812: data_o = 32'h00000000 /* 0xf710 */;
                15813: data_o = 32'h00000000 /* 0xf714 */;
                15814: data_o = 32'h00000000 /* 0xf718 */;
                15815: data_o = 32'h00000000 /* 0xf71c */;
                15816: data_o = 32'h00000000 /* 0xf720 */;
                15817: data_o = 32'h00000000 /* 0xf724 */;
                15818: data_o = 32'h00000000 /* 0xf728 */;
                15819: data_o = 32'h00000000 /* 0xf72c */;
                15820: data_o = 32'h00000000 /* 0xf730 */;
                15821: data_o = 32'h00000000 /* 0xf734 */;
                15822: data_o = 32'h00000000 /* 0xf738 */;
                15823: data_o = 32'h00000000 /* 0xf73c */;
                15824: data_o = 32'h00000000 /* 0xf740 */;
                15825: data_o = 32'h00000000 /* 0xf744 */;
                15826: data_o = 32'h00000000 /* 0xf748 */;
                15827: data_o = 32'h00000000 /* 0xf74c */;
                15828: data_o = 32'h00000000 /* 0xf750 */;
                15829: data_o = 32'h00000000 /* 0xf754 */;
                15830: data_o = 32'h00000000 /* 0xf758 */;
                15831: data_o = 32'h00000000 /* 0xf75c */;
                15832: data_o = 32'h00000000 /* 0xf760 */;
                15833: data_o = 32'h00000000 /* 0xf764 */;
                15834: data_o = 32'h00000000 /* 0xf768 */;
                15835: data_o = 32'h00000000 /* 0xf76c */;
                15836: data_o = 32'h00000000 /* 0xf770 */;
                15837: data_o = 32'h00000000 /* 0xf774 */;
                15838: data_o = 32'h00000000 /* 0xf778 */;
                15839: data_o = 32'h00000000 /* 0xf77c */;
                15840: data_o = 32'h00000000 /* 0xf780 */;
                15841: data_o = 32'h00000000 /* 0xf784 */;
                15842: data_o = 32'h00000000 /* 0xf788 */;
                15843: data_o = 32'h00000000 /* 0xf78c */;
                15844: data_o = 32'h00000000 /* 0xf790 */;
                15845: data_o = 32'h00000000 /* 0xf794 */;
                15846: data_o = 32'h00000000 /* 0xf798 */;
                15847: data_o = 32'h00000000 /* 0xf79c */;
                15848: data_o = 32'h00000000 /* 0xf7a0 */;
                15849: data_o = 32'h00000000 /* 0xf7a4 */;
                15850: data_o = 32'h00000000 /* 0xf7a8 */;
                15851: data_o = 32'h00000000 /* 0xf7ac */;
                15852: data_o = 32'h00000000 /* 0xf7b0 */;
                15853: data_o = 32'h00000000 /* 0xf7b4 */;
                15854: data_o = 32'h00000000 /* 0xf7b8 */;
                15855: data_o = 32'h00000000 /* 0xf7bc */;
                15856: data_o = 32'h00000000 /* 0xf7c0 */;
                15857: data_o = 32'h00000000 /* 0xf7c4 */;
                15858: data_o = 32'h00000000 /* 0xf7c8 */;
                15859: data_o = 32'h00000000 /* 0xf7cc */;
                15860: data_o = 32'h00000000 /* 0xf7d0 */;
                15861: data_o = 32'h00000000 /* 0xf7d4 */;
                15862: data_o = 32'h00000000 /* 0xf7d8 */;
                15863: data_o = 32'h00000000 /* 0xf7dc */;
                15864: data_o = 32'h00000000 /* 0xf7e0 */;
                15865: data_o = 32'h00000000 /* 0xf7e4 */;
                15866: data_o = 32'h00000000 /* 0xf7e8 */;
                15867: data_o = 32'h00000000 /* 0xf7ec */;
                15868: data_o = 32'h00000000 /* 0xf7f0 */;
                15869: data_o = 32'h00000000 /* 0xf7f4 */;
                15870: data_o = 32'h00000000 /* 0xf7f8 */;
                15871: data_o = 32'h00000000 /* 0xf7fc */;
                15872: data_o = 32'h00000000 /* 0xf800 */;
                15873: data_o = 32'h00000000 /* 0xf804 */;
                15874: data_o = 32'h00000000 /* 0xf808 */;
                15875: data_o = 32'h00000000 /* 0xf80c */;
                15876: data_o = 32'h00000000 /* 0xf810 */;
                15877: data_o = 32'h00000000 /* 0xf814 */;
                15878: data_o = 32'h00000000 /* 0xf818 */;
                15879: data_o = 32'h00000000 /* 0xf81c */;
                15880: data_o = 32'h00000000 /* 0xf820 */;
                15881: data_o = 32'h00000000 /* 0xf824 */;
                15882: data_o = 32'h00000000 /* 0xf828 */;
                15883: data_o = 32'h00000000 /* 0xf82c */;
                15884: data_o = 32'h00000000 /* 0xf830 */;
                15885: data_o = 32'h00000000 /* 0xf834 */;
                15886: data_o = 32'h00000000 /* 0xf838 */;
                15887: data_o = 32'h00000000 /* 0xf83c */;
                15888: data_o = 32'h00000000 /* 0xf840 */;
                15889: data_o = 32'h00000000 /* 0xf844 */;
                15890: data_o = 32'h00000000 /* 0xf848 */;
                15891: data_o = 32'h00000000 /* 0xf84c */;
                15892: data_o = 32'h00000000 /* 0xf850 */;
                15893: data_o = 32'h00000000 /* 0xf854 */;
                15894: data_o = 32'h00000000 /* 0xf858 */;
                15895: data_o = 32'h00000000 /* 0xf85c */;
                15896: data_o = 32'h00000000 /* 0xf860 */;
                15897: data_o = 32'h00000000 /* 0xf864 */;
                15898: data_o = 32'h00000000 /* 0xf868 */;
                15899: data_o = 32'h00000000 /* 0xf86c */;
                15900: data_o = 32'h00000000 /* 0xf870 */;
                15901: data_o = 32'h00000000 /* 0xf874 */;
                15902: data_o = 32'h00000000 /* 0xf878 */;
                15903: data_o = 32'h00000000 /* 0xf87c */;
                15904: data_o = 32'h00000000 /* 0xf880 */;
                15905: data_o = 32'h00000000 /* 0xf884 */;
                15906: data_o = 32'h00000000 /* 0xf888 */;
                15907: data_o = 32'h00000000 /* 0xf88c */;
                15908: data_o = 32'h00000000 /* 0xf890 */;
                15909: data_o = 32'h00000000 /* 0xf894 */;
                15910: data_o = 32'h00000000 /* 0xf898 */;
                15911: data_o = 32'h00000000 /* 0xf89c */;
                15912: data_o = 32'h00000000 /* 0xf8a0 */;
                15913: data_o = 32'h00000000 /* 0xf8a4 */;
                15914: data_o = 32'h00000000 /* 0xf8a8 */;
                15915: data_o = 32'h00000000 /* 0xf8ac */;
                15916: data_o = 32'h00000000 /* 0xf8b0 */;
                15917: data_o = 32'h00000000 /* 0xf8b4 */;
                15918: data_o = 32'h00000000 /* 0xf8b8 */;
                15919: data_o = 32'h00000000 /* 0xf8bc */;
                15920: data_o = 32'h00000000 /* 0xf8c0 */;
                15921: data_o = 32'h00000000 /* 0xf8c4 */;
                15922: data_o = 32'h00000000 /* 0xf8c8 */;
                15923: data_o = 32'h00000000 /* 0xf8cc */;
                15924: data_o = 32'h00000000 /* 0xf8d0 */;
                15925: data_o = 32'h00000000 /* 0xf8d4 */;
                15926: data_o = 32'h00000000 /* 0xf8d8 */;
                15927: data_o = 32'h00000000 /* 0xf8dc */;
                15928: data_o = 32'h00000000 /* 0xf8e0 */;
                15929: data_o = 32'h00000000 /* 0xf8e4 */;
                15930: data_o = 32'h00000000 /* 0xf8e8 */;
                15931: data_o = 32'h00000000 /* 0xf8ec */;
                15932: data_o = 32'h00000000 /* 0xf8f0 */;
                15933: data_o = 32'h00000000 /* 0xf8f4 */;
                15934: data_o = 32'h00000000 /* 0xf8f8 */;
                15935: data_o = 32'h00000000 /* 0xf8fc */;
                15936: data_o = 32'h00000000 /* 0xf900 */;
                15937: data_o = 32'h00000000 /* 0xf904 */;
                15938: data_o = 32'h00000000 /* 0xf908 */;
                15939: data_o = 32'h00000000 /* 0xf90c */;
                15940: data_o = 32'h00000000 /* 0xf910 */;
                15941: data_o = 32'h00000000 /* 0xf914 */;
                15942: data_o = 32'h00000000 /* 0xf918 */;
                15943: data_o = 32'h00000000 /* 0xf91c */;
                15944: data_o = 32'h00000000 /* 0xf920 */;
                15945: data_o = 32'h00000000 /* 0xf924 */;
                15946: data_o = 32'h00000000 /* 0xf928 */;
                15947: data_o = 32'h00000000 /* 0xf92c */;
                15948: data_o = 32'h00000000 /* 0xf930 */;
                15949: data_o = 32'h00000000 /* 0xf934 */;
                15950: data_o = 32'h00000000 /* 0xf938 */;
                15951: data_o = 32'h00000000 /* 0xf93c */;
                15952: data_o = 32'h00000000 /* 0xf940 */;
                15953: data_o = 32'h00000000 /* 0xf944 */;
                15954: data_o = 32'h00000000 /* 0xf948 */;
                15955: data_o = 32'h00000000 /* 0xf94c */;
                15956: data_o = 32'h00000000 /* 0xf950 */;
                15957: data_o = 32'h00000000 /* 0xf954 */;
                15958: data_o = 32'h00000000 /* 0xf958 */;
                15959: data_o = 32'h00000000 /* 0xf95c */;
                15960: data_o = 32'h00000000 /* 0xf960 */;
                15961: data_o = 32'h00000000 /* 0xf964 */;
                15962: data_o = 32'h00000000 /* 0xf968 */;
                15963: data_o = 32'h00000000 /* 0xf96c */;
                15964: data_o = 32'h00000000 /* 0xf970 */;
                15965: data_o = 32'h00000000 /* 0xf974 */;
                15966: data_o = 32'h00000000 /* 0xf978 */;
                15967: data_o = 32'h00000000 /* 0xf97c */;
                15968: data_o = 32'h00000000 /* 0xf980 */;
                15969: data_o = 32'h00000000 /* 0xf984 */;
                15970: data_o = 32'h00000000 /* 0xf988 */;
                15971: data_o = 32'h00000000 /* 0xf98c */;
                15972: data_o = 32'h00000000 /* 0xf990 */;
                15973: data_o = 32'h00000000 /* 0xf994 */;
                15974: data_o = 32'h00000000 /* 0xf998 */;
                15975: data_o = 32'h00000000 /* 0xf99c */;
                15976: data_o = 32'h00000000 /* 0xf9a0 */;
                15977: data_o = 32'h00000000 /* 0xf9a4 */;
                15978: data_o = 32'h00000000 /* 0xf9a8 */;
                15979: data_o = 32'h00000000 /* 0xf9ac */;
                15980: data_o = 32'h00000000 /* 0xf9b0 */;
                15981: data_o = 32'h00000000 /* 0xf9b4 */;
                15982: data_o = 32'h00000000 /* 0xf9b8 */;
                15983: data_o = 32'h00000000 /* 0xf9bc */;
                15984: data_o = 32'h00000000 /* 0xf9c0 */;
                15985: data_o = 32'h00000000 /* 0xf9c4 */;
                15986: data_o = 32'h00000000 /* 0xf9c8 */;
                15987: data_o = 32'h00000000 /* 0xf9cc */;
                15988: data_o = 32'h00000000 /* 0xf9d0 */;
                15989: data_o = 32'h00000000 /* 0xf9d4 */;
                15990: data_o = 32'h00000000 /* 0xf9d8 */;
                15991: data_o = 32'h00000000 /* 0xf9dc */;
                15992: data_o = 32'h00000000 /* 0xf9e0 */;
                15993: data_o = 32'h00000000 /* 0xf9e4 */;
                15994: data_o = 32'h00000000 /* 0xf9e8 */;
                15995: data_o = 32'h00000000 /* 0xf9ec */;
                15996: data_o = 32'h00000000 /* 0xf9f0 */;
                15997: data_o = 32'h00000000 /* 0xf9f4 */;
                15998: data_o = 32'h00000000 /* 0xf9f8 */;
                15999: data_o = 32'h00000000 /* 0xf9fc */;
                16000: data_o = 32'h00000000 /* 0xfa00 */;
                16001: data_o = 32'h00000000 /* 0xfa04 */;
                16002: data_o = 32'h00000000 /* 0xfa08 */;
                16003: data_o = 32'h00000000 /* 0xfa0c */;
                16004: data_o = 32'h00000000 /* 0xfa10 */;
                16005: data_o = 32'h00000000 /* 0xfa14 */;
                16006: data_o = 32'h00000000 /* 0xfa18 */;
                16007: data_o = 32'h00000000 /* 0xfa1c */;
                16008: data_o = 32'h00000000 /* 0xfa20 */;
                16009: data_o = 32'h00000000 /* 0xfa24 */;
                16010: data_o = 32'h00000000 /* 0xfa28 */;
                16011: data_o = 32'h00000000 /* 0xfa2c */;
                16012: data_o = 32'h00000000 /* 0xfa30 */;
                16013: data_o = 32'h00000000 /* 0xfa34 */;
                16014: data_o = 32'h00000000 /* 0xfa38 */;
                16015: data_o = 32'h00000000 /* 0xfa3c */;
                16016: data_o = 32'h00000000 /* 0xfa40 */;
                16017: data_o = 32'h00000000 /* 0xfa44 */;
                16018: data_o = 32'h00000000 /* 0xfa48 */;
                16019: data_o = 32'h00000000 /* 0xfa4c */;
                16020: data_o = 32'h00000000 /* 0xfa50 */;
                16021: data_o = 32'h00000000 /* 0xfa54 */;
                16022: data_o = 32'h00000000 /* 0xfa58 */;
                16023: data_o = 32'h00000000 /* 0xfa5c */;
                16024: data_o = 32'h00000000 /* 0xfa60 */;
                16025: data_o = 32'h00000000 /* 0xfa64 */;
                16026: data_o = 32'h00000000 /* 0xfa68 */;
                16027: data_o = 32'h00000000 /* 0xfa6c */;
                16028: data_o = 32'h00000000 /* 0xfa70 */;
                16029: data_o = 32'h00000000 /* 0xfa74 */;
                16030: data_o = 32'h00000000 /* 0xfa78 */;
                16031: data_o = 32'h00000000 /* 0xfa7c */;
                16032: data_o = 32'h00000000 /* 0xfa80 */;
                16033: data_o = 32'h00000000 /* 0xfa84 */;
                16034: data_o = 32'h00000000 /* 0xfa88 */;
                16035: data_o = 32'h00000000 /* 0xfa8c */;
                16036: data_o = 32'h00000000 /* 0xfa90 */;
                16037: data_o = 32'h00000000 /* 0xfa94 */;
                16038: data_o = 32'h00000000 /* 0xfa98 */;
                16039: data_o = 32'h00000000 /* 0xfa9c */;
                16040: data_o = 32'h00000000 /* 0xfaa0 */;
                16041: data_o = 32'h00000000 /* 0xfaa4 */;
                16042: data_o = 32'h00000000 /* 0xfaa8 */;
                16043: data_o = 32'h00000000 /* 0xfaac */;
                16044: data_o = 32'h00000000 /* 0xfab0 */;
                16045: data_o = 32'h00000000 /* 0xfab4 */;
                16046: data_o = 32'h00000000 /* 0xfab8 */;
                16047: data_o = 32'h00000000 /* 0xfabc */;
                16048: data_o = 32'h00000000 /* 0xfac0 */;
                16049: data_o = 32'h00000000 /* 0xfac4 */;
                16050: data_o = 32'h00000000 /* 0xfac8 */;
                16051: data_o = 32'h00000000 /* 0xfacc */;
                16052: data_o = 32'h00000000 /* 0xfad0 */;
                16053: data_o = 32'h00000000 /* 0xfad4 */;
                16054: data_o = 32'h00000000 /* 0xfad8 */;
                16055: data_o = 32'h00000000 /* 0xfadc */;
                16056: data_o = 32'h00000000 /* 0xfae0 */;
                16057: data_o = 32'h00000000 /* 0xfae4 */;
                16058: data_o = 32'h00000000 /* 0xfae8 */;
                16059: data_o = 32'h00000000 /* 0xfaec */;
                16060: data_o = 32'h00000000 /* 0xfaf0 */;
                16061: data_o = 32'h00000000 /* 0xfaf4 */;
                16062: data_o = 32'h00000000 /* 0xfaf8 */;
                16063: data_o = 32'h00000000 /* 0xfafc */;
                16064: data_o = 32'h00000000 /* 0xfb00 */;
                16065: data_o = 32'h00000000 /* 0xfb04 */;
                16066: data_o = 32'h00000000 /* 0xfb08 */;
                16067: data_o = 32'h00000000 /* 0xfb0c */;
                16068: data_o = 32'h00000000 /* 0xfb10 */;
                16069: data_o = 32'h00000000 /* 0xfb14 */;
                16070: data_o = 32'h00000000 /* 0xfb18 */;
                16071: data_o = 32'h00000000 /* 0xfb1c */;
                16072: data_o = 32'h00000000 /* 0xfb20 */;
                16073: data_o = 32'h00000000 /* 0xfb24 */;
                16074: data_o = 32'h00000000 /* 0xfb28 */;
                16075: data_o = 32'h00000000 /* 0xfb2c */;
                16076: data_o = 32'h00000000 /* 0xfb30 */;
                16077: data_o = 32'h00000000 /* 0xfb34 */;
                16078: data_o = 32'h00000000 /* 0xfb38 */;
                16079: data_o = 32'h00000000 /* 0xfb3c */;
                16080: data_o = 32'h00000000 /* 0xfb40 */;
                16081: data_o = 32'h00000000 /* 0xfb44 */;
                16082: data_o = 32'h00000000 /* 0xfb48 */;
                16083: data_o = 32'h00000000 /* 0xfb4c */;
                16084: data_o = 32'h00000000 /* 0xfb50 */;
                16085: data_o = 32'h00000000 /* 0xfb54 */;
                16086: data_o = 32'h00000000 /* 0xfb58 */;
                16087: data_o = 32'h00000000 /* 0xfb5c */;
                16088: data_o = 32'h00000000 /* 0xfb60 */;
                16089: data_o = 32'h00000000 /* 0xfb64 */;
                16090: data_o = 32'h00000000 /* 0xfb68 */;
                16091: data_o = 32'h00000000 /* 0xfb6c */;
                16092: data_o = 32'h00000000 /* 0xfb70 */;
                16093: data_o = 32'h00000000 /* 0xfb74 */;
                16094: data_o = 32'h00000000 /* 0xfb78 */;
                16095: data_o = 32'h00000000 /* 0xfb7c */;
                16096: data_o = 32'h00000000 /* 0xfb80 */;
                16097: data_o = 32'h00000000 /* 0xfb84 */;
                16098: data_o = 32'h00000000 /* 0xfb88 */;
                16099: data_o = 32'h00000000 /* 0xfb8c */;
                16100: data_o = 32'h00000000 /* 0xfb90 */;
                16101: data_o = 32'h00000000 /* 0xfb94 */;
                16102: data_o = 32'h00000000 /* 0xfb98 */;
                16103: data_o = 32'h00000000 /* 0xfb9c */;
                16104: data_o = 32'h00000000 /* 0xfba0 */;
                16105: data_o = 32'h00000000 /* 0xfba4 */;
                16106: data_o = 32'h00000000 /* 0xfba8 */;
                16107: data_o = 32'h00000000 /* 0xfbac */;
                16108: data_o = 32'h00000000 /* 0xfbb0 */;
                16109: data_o = 32'h00000000 /* 0xfbb4 */;
                16110: data_o = 32'h00000000 /* 0xfbb8 */;
                16111: data_o = 32'h00000000 /* 0xfbbc */;
                16112: data_o = 32'h00000000 /* 0xfbc0 */;
                16113: data_o = 32'h00000000 /* 0xfbc4 */;
                16114: data_o = 32'h00000000 /* 0xfbc8 */;
                16115: data_o = 32'h00000000 /* 0xfbcc */;
                16116: data_o = 32'h00000000 /* 0xfbd0 */;
                16117: data_o = 32'h00000000 /* 0xfbd4 */;
                16118: data_o = 32'h00000000 /* 0xfbd8 */;
                16119: data_o = 32'h00000000 /* 0xfbdc */;
                16120: data_o = 32'h00000000 /* 0xfbe0 */;
                16121: data_o = 32'h00000000 /* 0xfbe4 */;
                16122: data_o = 32'h00000000 /* 0xfbe8 */;
                16123: data_o = 32'h00000000 /* 0xfbec */;
                16124: data_o = 32'h00000000 /* 0xfbf0 */;
                16125: data_o = 32'h00000000 /* 0xfbf4 */;
                16126: data_o = 32'h00000000 /* 0xfbf8 */;
                16127: data_o = 32'h00000000 /* 0xfbfc */;
                16128: data_o = 32'h00000000 /* 0xfc00 */;
                16129: data_o = 32'h00000000 /* 0xfc04 */;
                16130: data_o = 32'h00000000 /* 0xfc08 */;
                16131: data_o = 32'h00000000 /* 0xfc0c */;
                16132: data_o = 32'h00000000 /* 0xfc10 */;
                16133: data_o = 32'h00000000 /* 0xfc14 */;
                16134: data_o = 32'h00000000 /* 0xfc18 */;
                16135: data_o = 32'h00000000 /* 0xfc1c */;
                16136: data_o = 32'h00000000 /* 0xfc20 */;
                16137: data_o = 32'h00000000 /* 0xfc24 */;
                16138: data_o = 32'h00000000 /* 0xfc28 */;
                16139: data_o = 32'h00000000 /* 0xfc2c */;
                16140: data_o = 32'h00000000 /* 0xfc30 */;
                16141: data_o = 32'h00000000 /* 0xfc34 */;
                16142: data_o = 32'h00000000 /* 0xfc38 */;
                16143: data_o = 32'h00000000 /* 0xfc3c */;
                16144: data_o = 32'h00000000 /* 0xfc40 */;
                16145: data_o = 32'h00000000 /* 0xfc44 */;
                16146: data_o = 32'h00000000 /* 0xfc48 */;
                16147: data_o = 32'h00000000 /* 0xfc4c */;
                16148: data_o = 32'h00000000 /* 0xfc50 */;
                16149: data_o = 32'h00000000 /* 0xfc54 */;
                16150: data_o = 32'h00000000 /* 0xfc58 */;
                16151: data_o = 32'h00000000 /* 0xfc5c */;
                16152: data_o = 32'h00000000 /* 0xfc60 */;
                16153: data_o = 32'h00000000 /* 0xfc64 */;
                16154: data_o = 32'h00000000 /* 0xfc68 */;
                16155: data_o = 32'h00000000 /* 0xfc6c */;
                16156: data_o = 32'h00000000 /* 0xfc70 */;
                16157: data_o = 32'h00000000 /* 0xfc74 */;
                16158: data_o = 32'h00000000 /* 0xfc78 */;
                16159: data_o = 32'h00000000 /* 0xfc7c */;
                16160: data_o = 32'h00000000 /* 0xfc80 */;
                16161: data_o = 32'h00000000 /* 0xfc84 */;
                16162: data_o = 32'h00000000 /* 0xfc88 */;
                16163: data_o = 32'h00000000 /* 0xfc8c */;
                16164: data_o = 32'h00000000 /* 0xfc90 */;
                16165: data_o = 32'h00000000 /* 0xfc94 */;
                16166: data_o = 32'h00000000 /* 0xfc98 */;
                16167: data_o = 32'h00000000 /* 0xfc9c */;
                16168: data_o = 32'h00000000 /* 0xfca0 */;
                16169: data_o = 32'h00000000 /* 0xfca4 */;
                16170: data_o = 32'h00000000 /* 0xfca8 */;
                16171: data_o = 32'h00000000 /* 0xfcac */;
                16172: data_o = 32'h00000000 /* 0xfcb0 */;
                16173: data_o = 32'h00000000 /* 0xfcb4 */;
                16174: data_o = 32'h00000000 /* 0xfcb8 */;
                16175: data_o = 32'h00000000 /* 0xfcbc */;
                16176: data_o = 32'h00000000 /* 0xfcc0 */;
                16177: data_o = 32'h00000000 /* 0xfcc4 */;
                16178: data_o = 32'h00000000 /* 0xfcc8 */;
                16179: data_o = 32'h00000000 /* 0xfccc */;
                16180: data_o = 32'h00000000 /* 0xfcd0 */;
                16181: data_o = 32'h00000000 /* 0xfcd4 */;
                16182: data_o = 32'h00000000 /* 0xfcd8 */;
                16183: data_o = 32'h00000000 /* 0xfcdc */;
                16184: data_o = 32'h00000000 /* 0xfce0 */;
                16185: data_o = 32'h00000000 /* 0xfce4 */;
                16186: data_o = 32'h00000000 /* 0xfce8 */;
                16187: data_o = 32'h00000000 /* 0xfcec */;
                16188: data_o = 32'h00000000 /* 0xfcf0 */;
                16189: data_o = 32'h00000000 /* 0xfcf4 */;
                16190: data_o = 32'h00000000 /* 0xfcf8 */;
                16191: data_o = 32'h00000000 /* 0xfcfc */;
                16192: data_o = 32'h00000000 /* 0xfd00 */;
                16193: data_o = 32'h00000000 /* 0xfd04 */;
                16194: data_o = 32'h00000000 /* 0xfd08 */;
                16195: data_o = 32'h00000000 /* 0xfd0c */;
                16196: data_o = 32'h00000000 /* 0xfd10 */;
                16197: data_o = 32'h00000000 /* 0xfd14 */;
                16198: data_o = 32'h00000000 /* 0xfd18 */;
                16199: data_o = 32'h00000000 /* 0xfd1c */;
                16200: data_o = 32'h00000000 /* 0xfd20 */;
                16201: data_o = 32'h00000000 /* 0xfd24 */;
                16202: data_o = 32'h00000000 /* 0xfd28 */;
                16203: data_o = 32'h00000000 /* 0xfd2c */;
                16204: data_o = 32'h00000000 /* 0xfd30 */;
                16205: data_o = 32'h00000000 /* 0xfd34 */;
                16206: data_o = 32'h00000000 /* 0xfd38 */;
                16207: data_o = 32'h00000000 /* 0xfd3c */;
                16208: data_o = 32'h00000000 /* 0xfd40 */;
                16209: data_o = 32'h00000000 /* 0xfd44 */;
                16210: data_o = 32'h00000000 /* 0xfd48 */;
                16211: data_o = 32'h00000000 /* 0xfd4c */;
                16212: data_o = 32'h00000000 /* 0xfd50 */;
                16213: data_o = 32'h00000000 /* 0xfd54 */;
                16214: data_o = 32'h00000000 /* 0xfd58 */;
                16215: data_o = 32'h00000000 /* 0xfd5c */;
                16216: data_o = 32'h00000000 /* 0xfd60 */;
                16217: data_o = 32'h00000000 /* 0xfd64 */;
                16218: data_o = 32'h00000000 /* 0xfd68 */;
                16219: data_o = 32'h00000000 /* 0xfd6c */;
                16220: data_o = 32'h00000000 /* 0xfd70 */;
                16221: data_o = 32'h00000000 /* 0xfd74 */;
                16222: data_o = 32'h00000000 /* 0xfd78 */;
                16223: data_o = 32'h00000000 /* 0xfd7c */;
                16224: data_o = 32'h00000000 /* 0xfd80 */;
                16225: data_o = 32'h00000000 /* 0xfd84 */;
                16226: data_o = 32'h00000000 /* 0xfd88 */;
                16227: data_o = 32'h00000000 /* 0xfd8c */;
                16228: data_o = 32'h00000000 /* 0xfd90 */;
                16229: data_o = 32'h00000000 /* 0xfd94 */;
                16230: data_o = 32'h00000000 /* 0xfd98 */;
                16231: data_o = 32'h00000000 /* 0xfd9c */;
                16232: data_o = 32'h00000000 /* 0xfda0 */;
                16233: data_o = 32'h00000000 /* 0xfda4 */;
                16234: data_o = 32'h00000000 /* 0xfda8 */;
                16235: data_o = 32'h00000000 /* 0xfdac */;
                16236: data_o = 32'h00000000 /* 0xfdb0 */;
                16237: data_o = 32'h00000000 /* 0xfdb4 */;
                16238: data_o = 32'h00000000 /* 0xfdb8 */;
                16239: data_o = 32'h00000000 /* 0xfdbc */;
                16240: data_o = 32'h00000000 /* 0xfdc0 */;
                16241: data_o = 32'h00000000 /* 0xfdc4 */;
                16242: data_o = 32'h00000000 /* 0xfdc8 */;
                16243: data_o = 32'h00000000 /* 0xfdcc */;
                16244: data_o = 32'h00000000 /* 0xfdd0 */;
                16245: data_o = 32'h00000000 /* 0xfdd4 */;
                16246: data_o = 32'h00000000 /* 0xfdd8 */;
                16247: data_o = 32'h00000000 /* 0xfddc */;
                16248: data_o = 32'h00000000 /* 0xfde0 */;
                16249: data_o = 32'h00000000 /* 0xfde4 */;
                16250: data_o = 32'h00000000 /* 0xfde8 */;
                16251: data_o = 32'h00000000 /* 0xfdec */;
                16252: data_o = 32'h00000000 /* 0xfdf0 */;
                16253: data_o = 32'h00000000 /* 0xfdf4 */;
                16254: data_o = 32'h00000000 /* 0xfdf8 */;
                16255: data_o = 32'h00000000 /* 0xfdfc */;
                16256: data_o = 32'h00000000 /* 0xfe00 */;
                16257: data_o = 32'h00000000 /* 0xfe04 */;
                16258: data_o = 32'h00000000 /* 0xfe08 */;
                16259: data_o = 32'h00000000 /* 0xfe0c */;
                16260: data_o = 32'h00000000 /* 0xfe10 */;
                16261: data_o = 32'h00000000 /* 0xfe14 */;
                16262: data_o = 32'h00000000 /* 0xfe18 */;
                16263: data_o = 32'h00000000 /* 0xfe1c */;
                16264: data_o = 32'h00000000 /* 0xfe20 */;
                16265: data_o = 32'h00000000 /* 0xfe24 */;
                16266: data_o = 32'h00000000 /* 0xfe28 */;
                16267: data_o = 32'h00000000 /* 0xfe2c */;
                16268: data_o = 32'h00000000 /* 0xfe30 */;
                16269: data_o = 32'h00000000 /* 0xfe34 */;
                16270: data_o = 32'h00000000 /* 0xfe38 */;
                16271: data_o = 32'h00000000 /* 0xfe3c */;
                16272: data_o = 32'h00000000 /* 0xfe40 */;
                16273: data_o = 32'h00000000 /* 0xfe44 */;
                16274: data_o = 32'h00000000 /* 0xfe48 */;
                16275: data_o = 32'h00000000 /* 0xfe4c */;
                16276: data_o = 32'h00000000 /* 0xfe50 */;
                16277: data_o = 32'h00000000 /* 0xfe54 */;
                16278: data_o = 32'h00000000 /* 0xfe58 */;
                16279: data_o = 32'h00000000 /* 0xfe5c */;
                16280: data_o = 32'h00000000 /* 0xfe60 */;
                16281: data_o = 32'h00000000 /* 0xfe64 */;
                16282: data_o = 32'h00000000 /* 0xfe68 */;
                16283: data_o = 32'h00000000 /* 0xfe6c */;
                16284: data_o = 32'h00000000 /* 0xfe70 */;
                16285: data_o = 32'h00000000 /* 0xfe74 */;
                16286: data_o = 32'h00000000 /* 0xfe78 */;
                16287: data_o = 32'h00000000 /* 0xfe7c */;
                16288: data_o = 32'h00000000 /* 0xfe80 */;
                16289: data_o = 32'h00000000 /* 0xfe84 */;
                16290: data_o = 32'h00000000 /* 0xfe88 */;
                16291: data_o = 32'h00000000 /* 0xfe8c */;
                16292: data_o = 32'h00000000 /* 0xfe90 */;
                16293: data_o = 32'h00000000 /* 0xfe94 */;
                16294: data_o = 32'h00000000 /* 0xfe98 */;
                16295: data_o = 32'h00000000 /* 0xfe9c */;
                16296: data_o = 32'h00000000 /* 0xfea0 */;
                16297: data_o = 32'h00000000 /* 0xfea4 */;
                16298: data_o = 32'h00000000 /* 0xfea8 */;
                16299: data_o = 32'h00000000 /* 0xfeac */;
                16300: data_o = 32'h00000000 /* 0xfeb0 */;
                16301: data_o = 32'h00000000 /* 0xfeb4 */;
                16302: data_o = 32'h00000000 /* 0xfeb8 */;
                16303: data_o = 32'h00000000 /* 0xfebc */;
                16304: data_o = 32'h00000000 /* 0xfec0 */;
                16305: data_o = 32'h00000000 /* 0xfec4 */;
                16306: data_o = 32'h00000000 /* 0xfec8 */;
                16307: data_o = 32'h00000000 /* 0xfecc */;
                16308: data_o = 32'h00000000 /* 0xfed0 */;
                16309: data_o = 32'h00000000 /* 0xfed4 */;
                16310: data_o = 32'h00000000 /* 0xfed8 */;
                16311: data_o = 32'h00000000 /* 0xfedc */;
                16312: data_o = 32'h00000000 /* 0xfee0 */;
                16313: data_o = 32'h00000000 /* 0xfee4 */;
                16314: data_o = 32'h00000000 /* 0xfee8 */;
                16315: data_o = 32'h00000000 /* 0xfeec */;
                16316: data_o = 32'h00000000 /* 0xfef0 */;
                16317: data_o = 32'h00000000 /* 0xfef4 */;
                16318: data_o = 32'h00000000 /* 0xfef8 */;
                16319: data_o = 32'h00000000 /* 0xfefc */;
                16320: data_o = 32'h00000000 /* 0xff00 */;
                16321: data_o = 32'h00000000 /* 0xff04 */;
                16322: data_o = 32'h00000000 /* 0xff08 */;
                16323: data_o = 32'h00000000 /* 0xff0c */;
                16324: data_o = 32'h00000000 /* 0xff10 */;
                16325: data_o = 32'h00000000 /* 0xff14 */;
                16326: data_o = 32'h00000000 /* 0xff18 */;
                16327: data_o = 32'h00000000 /* 0xff1c */;
                16328: data_o = 32'h00000000 /* 0xff20 */;
                16329: data_o = 32'h00000000 /* 0xff24 */;
                16330: data_o = 32'h00000000 /* 0xff28 */;
                16331: data_o = 32'h00000000 /* 0xff2c */;
                16332: data_o = 32'h00000000 /* 0xff30 */;
                16333: data_o = 32'h00000000 /* 0xff34 */;
                16334: data_o = 32'h00000000 /* 0xff38 */;
                16335: data_o = 32'h00000000 /* 0xff3c */;
                16336: data_o = 32'h00000000 /* 0xff40 */;
                16337: data_o = 32'h00000000 /* 0xff44 */;
                16338: data_o = 32'h00000000 /* 0xff48 */;
                16339: data_o = 32'h00000000 /* 0xff4c */;
                16340: data_o = 32'h00000000 /* 0xff50 */;
                16341: data_o = 32'h00000000 /* 0xff54 */;
                16342: data_o = 32'h00000000 /* 0xff58 */;
                16343: data_o = 32'h00000000 /* 0xff5c */;
                16344: data_o = 32'h00000000 /* 0xff60 */;
                16345: data_o = 32'h00000000 /* 0xff64 */;
                16346: data_o = 32'h00000000 /* 0xff68 */;
                16347: data_o = 32'h00000000 /* 0xff6c */;
                16348: data_o = 32'h00000000 /* 0xff70 */;
                16349: data_o = 32'h00000000 /* 0xff74 */;
                16350: data_o = 32'h00000000 /* 0xff78 */;
                16351: data_o = 32'h00000000 /* 0xff7c */;
                16352: data_o = 32'h00000000 /* 0xff80 */;
                16353: data_o = 32'h00000000 /* 0xff84 */;
                16354: data_o = 32'h00000000 /* 0xff88 */;
                16355: data_o = 32'h00000000 /* 0xff8c */;
                16356: data_o = 32'h00000000 /* 0xff90 */;
                16357: data_o = 32'h00000000 /* 0xff94 */;
                16358: data_o = 32'h00000000 /* 0xff98 */;
                16359: data_o = 32'h00000000 /* 0xff9c */;
                16360: data_o = 32'h00000000 /* 0xffa0 */;
                16361: data_o = 32'h00000000 /* 0xffa4 */;
                16362: data_o = 32'h00000000 /* 0xffa8 */;
                16363: data_o = 32'h00000000 /* 0xffac */;
                16364: data_o = 32'h00000000 /* 0xffb0 */;
                16365: data_o = 32'h00000000 /* 0xffb4 */;
                16366: data_o = 32'h00000000 /* 0xffb8 */;
                16367: data_o = 32'h00000000 /* 0xffbc */;
                16368: data_o = 32'h00000000 /* 0xffc0 */;
                16369: data_o = 32'h00000000 /* 0xffc4 */;
                16370: data_o = 32'h00000000 /* 0xffc8 */;
                16371: data_o = 32'h00000000 /* 0xffcc */;
                16372: data_o = 32'h00000000 /* 0xffd0 */;
                16373: data_o = 32'h00000000 /* 0xffd4 */;
                16374: data_o = 32'h00000000 /* 0xffd8 */;
                16375: data_o = 32'h00000000 /* 0xffdc */;
                16376: data_o = 32'h00000000 /* 0xffe0 */;
                16377: data_o = 32'h00000000 /* 0xffe4 */;
                16378: data_o = 32'h00000000 /* 0xffe8 */;
                16379: data_o = 32'h00000000 /* 0xffec */;
                16380: data_o = 32'h00000000 /* 0xfff0 */;
                16381: data_o = 32'h00000000 /* 0xfff4 */;
                16382: data_o = 32'h00000000 /* 0xfff8 */;
                16383: data_o = 32'h00000000 /* 0xfffc */;
                default: data_o = '0;
            endcase
        end

    endmodule
