`ifndef CHESHIRE_SVH
`define CHESHIRE_SVH


`define CHESHIRE_BASE_ADDR 64'h00000000
`define CHESHIRE_SIZE      64'h18000000


`define CHESHIRE_BOOT_ROM_BASE_ADDR 64'h02000000
`define CHESHIRE_BOOT_ROM_SIZE      64'h00040000


`define CHESHIRE_CHESHIRE_REGS_BASE_ADDR 64'h03000000
`define CHESHIRE_CHESHIRE_REGS_SIZE      64'h0000005C

`define CHESHIRE_CHESHIRE_REGS_SCRATCH_0_REG_ADDR   64'h03000000
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_0_REG_OFFSET 64'h00000000
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_1_REG_ADDR   64'h03000004
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_1_REG_OFFSET 64'h00000004
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_2_REG_ADDR   64'h03000008
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_2_REG_OFFSET 64'h00000008
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_3_REG_ADDR   64'h0300000C
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_3_REG_OFFSET 64'h0000000C
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_4_REG_ADDR   64'h03000010
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_4_REG_OFFSET 64'h00000010
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_5_REG_ADDR   64'h03000014
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_5_REG_OFFSET 64'h00000014
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_6_REG_ADDR   64'h03000018
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_6_REG_OFFSET 64'h00000018
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_7_REG_ADDR   64'h0300001C
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_7_REG_OFFSET 64'h0000001C
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_8_REG_ADDR   64'h03000020
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_8_REG_OFFSET 64'h00000020
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_9_REG_ADDR   64'h03000024
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_9_REG_OFFSET 64'h00000024
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_10_REG_ADDR   64'h03000028
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_10_REG_OFFSET 64'h00000028
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_11_REG_ADDR   64'h0300002C
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_11_REG_OFFSET 64'h0000002C
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_12_REG_ADDR   64'h03000030
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_12_REG_OFFSET 64'h00000030
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_13_REG_ADDR   64'h03000034
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_13_REG_OFFSET 64'h00000034
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_14_REG_ADDR   64'h03000038
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_14_REG_OFFSET 64'h00000038
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_15_REG_ADDR   64'h0300003C
`define CHESHIRE_CHESHIRE_REGS_SCRATCH_15_REG_OFFSET 64'h0000003C

`define CHESHIRE_CHESHIRE_REGS_BOOT_MODE_REG_ADDR   64'h03000040
`define CHESHIRE_CHESHIRE_REGS_BOOT_MODE_REG_OFFSET 64'h00000040

`define CHESHIRE_CHESHIRE_REGS_RTC_FREQ_REG_ADDR   64'h03000044
`define CHESHIRE_CHESHIRE_REGS_RTC_FREQ_REG_OFFSET 64'h00000044

`define CHESHIRE_CHESHIRE_REGS_PLATFORM_ROM_REG_ADDR   64'h03000048
`define CHESHIRE_CHESHIRE_REGS_PLATFORM_ROM_REG_OFFSET 64'h00000048

`define CHESHIRE_CHESHIRE_REGS_NUM_INT_HARTS_REG_ADDR   64'h0300004C
`define CHESHIRE_CHESHIRE_REGS_NUM_INT_HARTS_REG_OFFSET 64'h0000004C

`define CHESHIRE_CHESHIRE_REGS_HW_FEATURES_REG_ADDR   64'h03000050
`define CHESHIRE_CHESHIRE_REGS_HW_FEATURES_REG_OFFSET 64'h00000050

`define CHESHIRE_CHESHIRE_REGS_LLC_SIZE_REG_ADDR   64'h03000054
`define CHESHIRE_CHESHIRE_REGS_LLC_SIZE_REG_OFFSET 64'h00000054

`define CHESHIRE_CHESHIRE_REGS_VGA_PARAMS_REG_ADDR   64'h03000058
`define CHESHIRE_CHESHIRE_REGS_VGA_PARAMS_REG_OFFSET 64'h00000058


`define CHESHIRE_SERIAL_LINK_BASE_ADDR 64'h03006000
`define CHESHIRE_SERIAL_LINK_SIZE      64'h00000050


`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_BASE_ADDR 64'h03006000
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_SIZE      64'h00000050

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CTRL_REG_ADDR   64'h03006000
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CTRL_REG_OFFSET 64'h00000000

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_ISOLATED_REG_ADDR   64'h03006004
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_ISOLATED_REG_OFFSET 64'h00000004

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_TX_PHY_CLK_DIV_0_REG_ADDR   64'h03006008
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_TX_PHY_CLK_DIV_0_REG_OFFSET 64'h00000008

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_TX_PHY_CLK_START_0_REG_ADDR   64'h0300600C
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_TX_PHY_CLK_START_0_REG_OFFSET 64'h0000000C

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_TX_PHY_CLK_END_0_REG_ADDR   64'h03006010
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_TX_PHY_CLK_END_0_REG_OFFSET 64'h00000010

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_EN_REG_ADDR   64'h03006014
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_EN_REG_OFFSET 64'h00000014

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_IN_CH_SEL_REG_ADDR   64'h03006018
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_IN_CH_SEL_REG_OFFSET 64'h00000018

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_0_REG_ADDR   64'h0300601C
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_0_REG_OFFSET 64'h0000001C

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_IN_DATA_REG_ADDR   64'h03006020
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_IN_DATA_REG_OFFSET 64'h00000020

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_0_REG_ADDR   64'h03006024
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_0_REG_OFFSET 64'h00000024

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_REG_ADDR   64'h03006028
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_REG_OFFSET 64'h00000028

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_CTRL_REG_ADDR   64'h0300602C
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_CTRL_REG_OFFSET 64'h0000002C

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_OUT_EN_REG_ADDR   64'h03006030
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_RAW_MODE_OUT_EN_REG_OFFSET 64'h00000030

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_FLOW_CONTROL_FIFO_CLEAR_REG_ADDR   64'h03006034
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_FLOW_CONTROL_FIFO_CLEAR_REG_OFFSET 64'h00000034

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_TX_CFG_REG_ADDR   64'h03006038
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_TX_CFG_REG_OFFSET 64'h00000038

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_0_REG_ADDR   64'h0300603C
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_0_REG_OFFSET 64'h0000003C

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_TX_CTRL_REG_ADDR   64'h03006040
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_TX_CTRL_REG_OFFSET 64'h00000040

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_RX_CFG_REG_ADDR   64'h03006044
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_RX_CFG_REG_OFFSET 64'h00000044

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_RX_CTRL_REG_ADDR   64'h03006048
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_RX_CTRL_REG_OFFSET 64'h00000048

`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_0_REG_ADDR   64'h0300604C
`define CHESHIRE_SERIAL_LINK_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_0_REG_OFFSET 64'h0000004C


`define CHESHIRE_LLC_SPM_CACHED_BASE_ADDR 64'h10000000
`define CHESHIRE_LLC_SPM_CACHED_SIZE      64'h04000000


`define CHESHIRE_LLC_SPM_UNCACHED_BASE_ADDR 64'h14000000
`define CHESHIRE_LLC_SPM_UNCACHED_SIZE      64'h04000000


`endif /* CHESHIRE_SVH */
