// Copyright 2022 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
// Florian Zaruba <zarubaf@iis.ee.ethz.ch>
// Stefan Mach <smach@iis.ee.ethz.ch>
// Thomas Benz <tbenz@iis.ee.ethz.ch>
// Paul Scheffler <paulsc@iis.ee.ethz.ch>
// Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
//
// AUTOMATICALLY GENERATED by gen_bootrom.py; edit the script instead.

module cheshire_bootrom #(
    parameter int unsigned AddrWidth = 32,
    parameter int unsigned DataWidth = 32
)(
    input  logic                 clk_i,
    input  logic                 rst_ni,
    input  logic                 req_i,
    input  logic [AddrWidth-1:0] addr_i,
    output logic [DataWidth-1:0] data_o
);
    localparam unsigned NumWords = 64;
    logic [$clog2(NumWords)-1:0] word;

    assign word = addr_i / (DataWidth / 8);

    always_comb begin
        data_o = '0;
        unique case (word)
        000: data_o = 32'h6f006117 /* 0x0000 */;
            001: data_o = 32'hff810113 /* 0x0004 */;
            002: data_o = 32'h00000197 /* 0x0008 */;
            003: data_o = 32'h0c818193 /* 0x000c */;
            004: data_o = 32'h42014081 /* 0x0010 */;
            005: data_o = 32'h43014281 /* 0x0014 */;
            006: data_o = 32'h44014381 /* 0x0018 */;
            007: data_o = 32'h45014481 /* 0x001c */;
            008: data_o = 32'h46014581 /* 0x0020 */;
            009: data_o = 32'h47014681 /* 0x0024 */;
            010: data_o = 32'h48014781 /* 0x0028 */;
            011: data_o = 32'h49014881 /* 0x002c */;
            012: data_o = 32'h4a014981 /* 0x0030 */;
            013: data_o = 32'h4b014a81 /* 0x0034 */;
            014: data_o = 32'h4c014b81 /* 0x0038 */;
            015: data_o = 32'h4d014c81 /* 0x003c */;
            016: data_o = 32'h4e014d81 /* 0x0040 */;
            017: data_o = 32'h4f014e81 /* 0x0044 */;
            018: data_o = 32'h12974f81 /* 0x0048 */;
            019: data_o = 32'h82930100 /* 0x004c */;
            020: data_o = 32'h537dfb62 /* 0x0050 */;
            021: data_o = 32'h0062a023 /* 0x0054 */;
            022: data_o = 32'h0062a223 /* 0x0058 */;
            023: data_o = 32'ha8234305 /* 0x005c */;
            024: data_o = 32'h42810062 /* 0x0060 */;
            025: data_o = 32'h100f4301 /* 0x0064 */;
            026: data_o = 32'h00ef0000 /* 0x0068 */;
            027: data_o = 32'ha00903c0 /* 0x006c */;
            028: data_o = 32'h65130506 /* 0x0070 */;
            029: data_o = 32'h02970015 /* 0x0074 */;
            030: data_o = 32'h82930100 /* 0x0078 */;
            031: data_o = 32'ha223f8a2 /* 0x007c */;
            032: data_o = 32'h007300a2 /* 0x0080 */;
            033: data_o = 32'hbff51050 /* 0x0084 */;
            034: data_o = 32'h020007b7 /* 0x0088 */;
            035: data_o = 32'h00078793 /* 0x008c */;
            036: data_o = 32'hdf7d4798 /* 0x0090 */;
            037: data_o = 32'h0ff0000f /* 0x0094 */;
            038: data_o = 32'h278143dc /* 0x0098 */;
            039: data_o = 32'h0000100f /* 0x009c */;
            040: data_o = 32'h93811782 /* 0x00a0 */;
            041: data_o = 32'h07b78782 /* 0x00a4 */;
            042: data_o = 32'h87930200 /* 0x00a8 */;
            043: data_o = 32'h4bd80007 /* 0x00ac */;
            044: data_o = 32'h079b579c /* 0x00b0 */;
            045: data_o = 32'h4709fff7 /* 0x00b4 */;
            046: data_o = 32'h00f77a63 /* 0x00b8 */;
            047: data_o = 32'he4061141 /* 0x00bc */;
            048: data_o = 32'hfc9ff0ef /* 0x00c0 */;
            049: data_o = 32'h250160a2 /* 0x00c4 */;
            050: data_o = 32'h80820141 /* 0x00c8 */;
            051: data_o = 32'h80824501 /* 0x00cc */;
            052: data_o = 32'h00000000 /* 0x00d0 */;
            053: data_o = 32'h00000000 /* 0x00d4 */;
            054: data_o = 32'h00000000 /* 0x00d8 */;
            055: data_o = 32'h00000000 /* 0x00dc */;
            056: data_o = 32'h00000000 /* 0x00e0 */;
            057: data_o = 32'h00000000 /* 0x00e4 */;
            058: data_o = 32'h00000000 /* 0x00e8 */;
            059: data_o = 32'h00000000 /* 0x00ec */;
            060: data_o = 32'h00000000 /* 0x00f0 */;
            061: data_o = 32'h00000000 /* 0x00f4 */;
            062: data_o = 32'h00000000 /* 0x00f8 */;
            063: data_o = 32'h00000000 /* 0x00fc */;
            default: data_o = '0;
        endcase
    end

endmodule
